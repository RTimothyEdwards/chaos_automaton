VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chaos_subarray
  CLASS BLOCK ;
  FOREIGN chaos_subarray ;
  ORIGIN 0.000 0.000 ;
  SIZE 825.000 BY 585.000 ;
  PIN hold
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END hold
  PIN iclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END iclk
  PIN idata
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END idata
  PIN ieast[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 13.640 825.000 14.240 ;
    END
  END ieast[0]
  PIN ieast[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 40.160 825.000 40.760 ;
    END
  END ieast[1]
  PIN ieast[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 66.680 825.000 67.280 ;
    END
  END ieast[2]
  PIN ieast[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 93.200 825.000 93.800 ;
    END
  END ieast[3]
  PIN ieast[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 119.720 825.000 120.320 ;
    END
  END ieast[4]
  PIN ieast[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 146.240 825.000 146.840 ;
    END
  END ieast[5]
  PIN ieast[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 172.760 825.000 173.360 ;
    END
  END ieast[6]
  PIN ieast[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 199.280 825.000 199.880 ;
    END
  END ieast[7]
  PIN ieast[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 225.800 825.000 226.400 ;
    END
  END ieast[8]
  PIN ieast[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 252.320 825.000 252.920 ;
    END
  END ieast[9]
  PIN inorth[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 581.000 801.230 585.000 ;
    END
  END inorth[0]
  PIN inorth[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 581.000 760.290 585.000 ;
    END
  END inorth[1]
  PIN inorth[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 581.000 719.350 585.000 ;
    END
  END inorth[2]
  PIN inorth[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 581.000 678.410 585.000 ;
    END
  END inorth[3]
  PIN inorth[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 581.000 637.470 585.000 ;
    END
  END inorth[4]
  PIN inorth[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 581.000 596.530 585.000 ;
    END
  END inorth[5]
  PIN inorth[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 581.000 555.590 585.000 ;
    END
  END inorth[6]
  PIN inorth[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 581.000 514.650 585.000 ;
    END
  END inorth[7]
  PIN inorth[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 581.000 473.710 585.000 ;
    END
  END inorth[8]
  PIN inorth[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 581.000 432.770 585.000 ;
    END
  END inorth[9]
  PIN isouth[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END isouth[0]
  PIN isouth[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END isouth[1]
  PIN isouth[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END isouth[2]
  PIN isouth[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END isouth[3]
  PIN isouth[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END isouth[4]
  PIN isouth[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END isouth[5]
  PIN isouth[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END isouth[6]
  PIN isouth[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END isouth[7]
  PIN isouth[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END isouth[8]
  PIN isouth[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END isouth[9]
  PIN iwest[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 570.560 4.000 571.160 ;
    END
  END iwest[0]
  PIN iwest[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END iwest[1]
  PIN iwest[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 517.520 4.000 518.120 ;
    END
  END iwest[2]
  PIN iwest[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END iwest[3]
  PIN iwest[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 464.480 4.000 465.080 ;
    END
  END iwest[4]
  PIN iwest[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END iwest[5]
  PIN iwest[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END iwest[6]
  PIN iwest[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END iwest[7]
  PIN iwest[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END iwest[8]
  PIN iwest[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END iwest[9]
  PIN oclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 544.040 825.000 544.640 ;
    END
  END oclk
  PIN odata
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 570.560 825.000 571.160 ;
    END
  END odata
  PIN oeast[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 278.840 825.000 279.440 ;
    END
  END oeast[0]
  PIN oeast[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 305.360 825.000 305.960 ;
    END
  END oeast[1]
  PIN oeast[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 331.880 825.000 332.480 ;
    END
  END oeast[2]
  PIN oeast[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 358.400 825.000 359.000 ;
    END
  END oeast[3]
  PIN oeast[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 384.920 825.000 385.520 ;
    END
  END oeast[4]
  PIN oeast[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 411.440 825.000 412.040 ;
    END
  END oeast[5]
  PIN oeast[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 437.960 825.000 438.560 ;
    END
  END oeast[6]
  PIN oeast[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 464.480 825.000 465.080 ;
    END
  END oeast[7]
  PIN oeast[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 491.000 825.000 491.600 ;
    END
  END oeast[8]
  PIN oeast[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.000 517.520 825.000 518.120 ;
    END
  END oeast[9]
  PIN onorth[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 581.000 391.830 585.000 ;
    END
  END onorth[0]
  PIN onorth[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 581.000 350.890 585.000 ;
    END
  END onorth[1]
  PIN onorth[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 581.000 309.950 585.000 ;
    END
  END onorth[2]
  PIN onorth[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 581.000 269.010 585.000 ;
    END
  END onorth[3]
  PIN onorth[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 581.000 228.070 585.000 ;
    END
  END onorth[4]
  PIN onorth[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 581.000 187.130 585.000 ;
    END
  END onorth[5]
  PIN onorth[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 581.000 146.190 585.000 ;
    END
  END onorth[6]
  PIN onorth[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 581.000 105.250 585.000 ;
    END
  END onorth[7]
  PIN onorth[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 581.000 64.310 585.000 ;
    END
  END onorth[8]
  PIN onorth[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 581.000 23.370 585.000 ;
    END
  END onorth[9]
  PIN osouth[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END osouth[0]
  PIN osouth[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END osouth[1]
  PIN osouth[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END osouth[2]
  PIN osouth[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END osouth[3]
  PIN osouth[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 0.000 617.230 4.000 ;
    END
  END osouth[4]
  PIN osouth[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END osouth[5]
  PIN osouth[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 0.000 691.750 4.000 ;
    END
  END osouth[6]
  PIN osouth[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 0.000 729.010 4.000 ;
    END
  END osouth[7]
  PIN osouth[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END osouth[8]
  PIN osouth[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.250 0.000 803.530 4.000 ;
    END
  END osouth[9]
  PIN owest[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END owest[0]
  PIN owest[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END owest[1]
  PIN owest[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END owest[2]
  PIN owest[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END owest[3]
  PIN owest[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END owest[4]
  PIN owest[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END owest[5]
  PIN owest[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END owest[6]
  PIN owest[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END owest[7]
  PIN owest[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END owest[8]
  PIN owest[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END owest[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.340 10.640 34.340 574.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 162.940 10.640 187.940 574.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.540 10.640 341.540 574.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 470.140 10.640 495.140 574.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.740 10.640 648.740 574.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 777.340 10.640 802.340 574.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 86.140 10.640 111.140 574.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 239.740 10.640 264.740 574.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 393.340 10.640 418.340 574.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.940 10.640 571.940 574.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 700.540 10.640 725.540 574.160 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 819.260 574.005 ;
      LAYER met1 ;
        RECT 2.830 8.880 819.260 575.920 ;
      LAYER met2 ;
        RECT 2.860 580.720 22.810 581.810 ;
        RECT 23.650 580.720 63.750 581.810 ;
        RECT 64.590 580.720 104.690 581.810 ;
        RECT 105.530 580.720 145.630 581.810 ;
        RECT 146.470 580.720 186.570 581.810 ;
        RECT 187.410 580.720 227.510 581.810 ;
        RECT 228.350 580.720 268.450 581.810 ;
        RECT 269.290 580.720 309.390 581.810 ;
        RECT 310.230 580.720 350.330 581.810 ;
        RECT 351.170 580.720 391.270 581.810 ;
        RECT 392.110 580.720 432.210 581.810 ;
        RECT 433.050 580.720 473.150 581.810 ;
        RECT 473.990 580.720 514.090 581.810 ;
        RECT 514.930 580.720 555.030 581.810 ;
        RECT 555.870 580.720 595.970 581.810 ;
        RECT 596.810 580.720 636.910 581.810 ;
        RECT 637.750 580.720 677.850 581.810 ;
        RECT 678.690 580.720 718.790 581.810 ;
        RECT 719.630 580.720 759.730 581.810 ;
        RECT 760.570 580.720 800.670 581.810 ;
        RECT 801.510 580.720 818.240 581.810 ;
        RECT 2.860 4.280 818.240 580.720 ;
        RECT 2.860 3.670 20.510 4.280 ;
        RECT 21.350 3.670 57.770 4.280 ;
        RECT 58.610 3.670 95.030 4.280 ;
        RECT 95.870 3.670 132.290 4.280 ;
        RECT 133.130 3.670 169.550 4.280 ;
        RECT 170.390 3.670 206.810 4.280 ;
        RECT 207.650 3.670 244.070 4.280 ;
        RECT 244.910 3.670 281.330 4.280 ;
        RECT 282.170 3.670 318.590 4.280 ;
        RECT 319.430 3.670 355.850 4.280 ;
        RECT 356.690 3.670 393.110 4.280 ;
        RECT 393.950 3.670 430.370 4.280 ;
        RECT 431.210 3.670 467.630 4.280 ;
        RECT 468.470 3.670 504.890 4.280 ;
        RECT 505.730 3.670 542.150 4.280 ;
        RECT 542.990 3.670 579.410 4.280 ;
        RECT 580.250 3.670 616.670 4.280 ;
        RECT 617.510 3.670 653.930 4.280 ;
        RECT 654.770 3.670 691.190 4.280 ;
        RECT 692.030 3.670 728.450 4.280 ;
        RECT 729.290 3.670 765.710 4.280 ;
        RECT 766.550 3.670 802.970 4.280 ;
        RECT 803.810 3.670 818.240 4.280 ;
      LAYER met3 ;
        RECT 4.000 571.560 821.000 574.085 ;
        RECT 4.400 570.160 820.600 571.560 ;
        RECT 4.000 545.040 821.000 570.160 ;
        RECT 4.400 543.640 820.600 545.040 ;
        RECT 4.000 518.520 821.000 543.640 ;
        RECT 4.400 517.120 820.600 518.520 ;
        RECT 4.000 492.000 821.000 517.120 ;
        RECT 4.400 490.600 820.600 492.000 ;
        RECT 4.000 465.480 821.000 490.600 ;
        RECT 4.400 464.080 820.600 465.480 ;
        RECT 4.000 438.960 821.000 464.080 ;
        RECT 4.400 437.560 820.600 438.960 ;
        RECT 4.000 412.440 821.000 437.560 ;
        RECT 4.400 411.040 820.600 412.440 ;
        RECT 4.000 385.920 821.000 411.040 ;
        RECT 4.400 384.520 820.600 385.920 ;
        RECT 4.000 359.400 821.000 384.520 ;
        RECT 4.400 358.000 820.600 359.400 ;
        RECT 4.000 332.880 821.000 358.000 ;
        RECT 4.400 331.480 820.600 332.880 ;
        RECT 4.000 306.360 821.000 331.480 ;
        RECT 4.400 304.960 820.600 306.360 ;
        RECT 4.000 279.840 821.000 304.960 ;
        RECT 4.400 278.440 820.600 279.840 ;
        RECT 4.000 253.320 821.000 278.440 ;
        RECT 4.400 251.920 820.600 253.320 ;
        RECT 4.000 226.800 821.000 251.920 ;
        RECT 4.400 225.400 820.600 226.800 ;
        RECT 4.000 200.280 821.000 225.400 ;
        RECT 4.400 198.880 820.600 200.280 ;
        RECT 4.000 173.760 821.000 198.880 ;
        RECT 4.400 172.360 820.600 173.760 ;
        RECT 4.000 147.240 821.000 172.360 ;
        RECT 4.400 145.840 820.600 147.240 ;
        RECT 4.000 120.720 821.000 145.840 ;
        RECT 4.400 119.320 820.600 120.720 ;
        RECT 4.000 94.200 821.000 119.320 ;
        RECT 4.400 92.800 820.600 94.200 ;
        RECT 4.000 67.680 821.000 92.800 ;
        RECT 4.400 66.280 820.600 67.680 ;
        RECT 4.000 41.160 821.000 66.280 ;
        RECT 4.400 39.760 820.600 41.160 ;
        RECT 4.000 14.640 821.000 39.760 ;
        RECT 4.400 13.240 820.600 14.640 ;
        RECT 4.000 10.715 821.000 13.240 ;
      LAYER met4 ;
        RECT 7.655 13.095 8.940 567.625 ;
        RECT 34.740 13.095 85.740 567.625 ;
        RECT 111.540 13.095 162.540 567.625 ;
        RECT 188.340 13.095 239.340 567.625 ;
        RECT 265.140 13.095 316.140 567.625 ;
        RECT 341.940 13.095 392.940 567.625 ;
        RECT 418.740 13.095 469.740 567.625 ;
        RECT 495.540 13.095 546.540 567.625 ;
        RECT 572.340 13.095 623.340 567.625 ;
        RECT 649.140 13.095 700.140 567.625 ;
        RECT 725.940 13.095 776.940 567.625 ;
        RECT 802.740 13.095 813.905 567.625 ;
  END
END chaos_subarray
END LIBRARY

