magic
tech sky130B
magscale 1 2
timestamp 1659731860
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 1640 178848 117552
<< metal2 >>
rect 5170 119200 5226 120000
rect 14094 119200 14150 120000
rect 23018 119200 23074 120000
rect 31942 119200 31998 120000
rect 40866 119200 40922 120000
rect 49790 119200 49846 120000
rect 58714 119200 58770 120000
rect 67638 119200 67694 120000
rect 76562 119200 76618 120000
rect 85486 119200 85542 120000
rect 94410 119200 94466 120000
rect 103334 119200 103390 120000
rect 112258 119200 112314 120000
rect 121182 119200 121238 120000
rect 130106 119200 130162 120000
rect 139030 119200 139086 120000
rect 147954 119200 148010 120000
rect 156878 119200 156934 120000
rect 165802 119200 165858 120000
rect 174726 119200 174782 120000
rect 4986 0 5042 800
rect 13082 0 13138 800
rect 21178 0 21234 800
rect 29274 0 29330 800
rect 37370 0 37426 800
rect 45466 0 45522 800
rect 53562 0 53618 800
rect 61658 0 61714 800
rect 69754 0 69810 800
rect 77850 0 77906 800
rect 85946 0 86002 800
rect 94042 0 94098 800
rect 102138 0 102194 800
rect 110234 0 110290 800
rect 118330 0 118386 800
rect 126426 0 126482 800
rect 134522 0 134578 800
rect 142618 0 142674 800
rect 150714 0 150770 800
rect 158810 0 158866 800
rect 166906 0 166962 800
rect 175002 0 175058 800
<< obsm2 >>
rect 1398 119144 5114 119354
rect 5282 119144 14038 119354
rect 14206 119144 22962 119354
rect 23130 119144 31886 119354
rect 32054 119144 40810 119354
rect 40978 119144 49734 119354
rect 49902 119144 58658 119354
rect 58826 119144 67582 119354
rect 67750 119144 76506 119354
rect 76674 119144 85430 119354
rect 85598 119144 94354 119354
rect 94522 119144 103278 119354
rect 103446 119144 112202 119354
rect 112370 119144 121126 119354
rect 121294 119144 130050 119354
rect 130218 119144 138974 119354
rect 139142 119144 147898 119354
rect 148066 119144 156822 119354
rect 156990 119144 165746 119354
rect 165914 119144 174670 119354
rect 174838 119144 178462 119354
rect 1398 856 178462 119144
rect 1398 800 4930 856
rect 5098 800 13026 856
rect 13194 800 21122 856
rect 21290 800 29218 856
rect 29386 800 37314 856
rect 37482 800 45410 856
rect 45578 800 53506 856
rect 53674 800 61602 856
rect 61770 800 69698 856
rect 69866 800 77794 856
rect 77962 800 85890 856
rect 86058 800 93986 856
rect 94154 800 102082 856
rect 102250 800 110178 856
rect 110346 800 118274 856
rect 118442 800 126370 856
rect 126538 800 134466 856
rect 134634 800 142562 856
rect 142730 800 150658 856
rect 150826 800 158754 856
rect 158922 800 166850 856
rect 167018 800 174946 856
rect 175114 800 178462 856
<< metal3 >>
rect 0 116968 800 117088
rect 179200 116968 180000 117088
rect 0 111528 800 111648
rect 179200 111528 180000 111648
rect 0 106088 800 106208
rect 179200 106088 180000 106208
rect 0 100648 800 100768
rect 179200 100648 180000 100768
rect 0 95208 800 95328
rect 179200 95208 180000 95328
rect 0 89768 800 89888
rect 179200 89768 180000 89888
rect 0 84328 800 84448
rect 179200 84328 180000 84448
rect 0 78888 800 79008
rect 179200 78888 180000 79008
rect 0 73448 800 73568
rect 179200 73448 180000 73568
rect 0 68008 800 68128
rect 179200 68008 180000 68128
rect 0 62568 800 62688
rect 179200 62568 180000 62688
rect 0 57128 800 57248
rect 179200 57128 180000 57248
rect 0 51688 800 51808
rect 179200 51688 180000 51808
rect 0 46248 800 46368
rect 179200 46248 180000 46368
rect 0 40808 800 40928
rect 179200 40808 180000 40928
rect 0 35368 800 35488
rect 179200 35368 180000 35488
rect 0 29928 800 30048
rect 179200 29928 180000 30048
rect 0 24488 800 24608
rect 179200 24488 180000 24608
rect 0 19048 800 19168
rect 179200 19048 180000 19168
rect 0 13608 800 13728
rect 179200 13608 180000 13728
rect 0 8168 800 8288
rect 179200 8168 180000 8288
rect 0 2728 800 2848
rect 179200 2728 180000 2848
<< obsm3 >>
rect 800 117168 179200 117537
rect 880 116888 179120 117168
rect 800 111728 179200 116888
rect 880 111448 179120 111728
rect 800 106288 179200 111448
rect 880 106008 179120 106288
rect 800 100848 179200 106008
rect 880 100568 179120 100848
rect 800 95408 179200 100568
rect 880 95128 179120 95408
rect 800 89968 179200 95128
rect 880 89688 179120 89968
rect 800 84528 179200 89688
rect 880 84248 179120 84528
rect 800 79088 179200 84248
rect 880 78808 179120 79088
rect 800 73648 179200 78808
rect 880 73368 179120 73648
rect 800 68208 179200 73368
rect 880 67928 179120 68208
rect 800 62768 179200 67928
rect 880 62488 179120 62768
rect 800 57328 179200 62488
rect 880 57048 179120 57328
rect 800 51888 179200 57048
rect 880 51608 179120 51888
rect 800 46448 179200 51608
rect 880 46168 179120 46448
rect 800 41008 179200 46168
rect 880 40728 179120 41008
rect 800 35568 179200 40728
rect 880 35288 179120 35568
rect 800 30128 179200 35288
rect 880 29848 179120 30128
rect 800 24688 179200 29848
rect 880 24408 179120 24688
rect 800 19248 179200 24408
rect 880 18968 179120 19248
rect 800 13808 179200 18968
rect 880 13528 179120 13808
rect 800 8368 179200 13528
rect 880 8088 179120 8368
rect 800 2928 179200 8088
rect 880 2648 179120 2928
rect 800 2143 179200 2648
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 2083 14043 4128 106317
rect 4608 14043 19488 106317
rect 19968 14043 34848 106317
rect 35328 14043 50208 106317
rect 50688 14043 65568 106317
rect 66048 14043 80928 106317
rect 81408 14043 96288 106317
rect 96768 14043 111648 106317
rect 112128 14043 127008 106317
rect 127488 14043 142368 106317
rect 142848 14043 157728 106317
rect 158208 14043 173088 106317
rect 173568 14043 177869 106317
<< metal5 >>
rect 1056 112572 178896 112892
rect 1056 97254 178896 97574
rect 1056 81936 178896 82256
rect 1056 66618 178896 66938
rect 1056 51300 178896 51620
rect 1056 35982 178896 36302
rect 1056 20664 178896 20984
rect 1056 5346 178896 5666
<< labels >>
rlabel metal2 s 4986 0 5042 800 6 hold
port 1 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 iclk
port 2 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 idata
port 3 nsew signal input
rlabel metal3 s 179200 2728 180000 2848 6 ieast[0]
port 4 nsew signal input
rlabel metal3 s 179200 8168 180000 8288 6 ieast[1]
port 5 nsew signal input
rlabel metal3 s 179200 13608 180000 13728 6 ieast[2]
port 6 nsew signal input
rlabel metal3 s 179200 19048 180000 19168 6 ieast[3]
port 7 nsew signal input
rlabel metal3 s 179200 24488 180000 24608 6 ieast[4]
port 8 nsew signal input
rlabel metal3 s 179200 29928 180000 30048 6 ieast[5]
port 9 nsew signal input
rlabel metal3 s 179200 35368 180000 35488 6 ieast[6]
port 10 nsew signal input
rlabel metal3 s 179200 40808 180000 40928 6 ieast[7]
port 11 nsew signal input
rlabel metal3 s 179200 46248 180000 46368 6 ieast[8]
port 12 nsew signal input
rlabel metal3 s 179200 51688 180000 51808 6 ieast[9]
port 13 nsew signal input
rlabel metal2 s 174726 119200 174782 120000 6 inorth[0]
port 14 nsew signal input
rlabel metal2 s 165802 119200 165858 120000 6 inorth[1]
port 15 nsew signal input
rlabel metal2 s 156878 119200 156934 120000 6 inorth[2]
port 16 nsew signal input
rlabel metal2 s 147954 119200 148010 120000 6 inorth[3]
port 17 nsew signal input
rlabel metal2 s 139030 119200 139086 120000 6 inorth[4]
port 18 nsew signal input
rlabel metal2 s 130106 119200 130162 120000 6 inorth[5]
port 19 nsew signal input
rlabel metal2 s 121182 119200 121238 120000 6 inorth[6]
port 20 nsew signal input
rlabel metal2 s 112258 119200 112314 120000 6 inorth[7]
port 21 nsew signal input
rlabel metal2 s 103334 119200 103390 120000 6 inorth[8]
port 22 nsew signal input
rlabel metal2 s 94410 119200 94466 120000 6 inorth[9]
port 23 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 isouth[0]
port 24 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 isouth[1]
port 25 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 isouth[2]
port 26 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 isouth[3]
port 27 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 isouth[4]
port 28 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 isouth[5]
port 29 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 isouth[6]
port 30 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 isouth[7]
port 31 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 isouth[8]
port 32 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 isouth[9]
port 33 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 iwest[0]
port 34 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 iwest[1]
port 35 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 iwest[2]
port 36 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 iwest[3]
port 37 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 iwest[4]
port 38 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 iwest[5]
port 39 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 iwest[6]
port 40 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 iwest[7]
port 41 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 iwest[8]
port 42 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 iwest[9]
port 43 nsew signal input
rlabel metal3 s 179200 111528 180000 111648 6 oclk
port 44 nsew signal output
rlabel metal3 s 179200 116968 180000 117088 6 odata
port 45 nsew signal output
rlabel metal3 s 179200 57128 180000 57248 6 oeast[0]
port 46 nsew signal output
rlabel metal3 s 179200 62568 180000 62688 6 oeast[1]
port 47 nsew signal output
rlabel metal3 s 179200 68008 180000 68128 6 oeast[2]
port 48 nsew signal output
rlabel metal3 s 179200 73448 180000 73568 6 oeast[3]
port 49 nsew signal output
rlabel metal3 s 179200 78888 180000 79008 6 oeast[4]
port 50 nsew signal output
rlabel metal3 s 179200 84328 180000 84448 6 oeast[5]
port 51 nsew signal output
rlabel metal3 s 179200 89768 180000 89888 6 oeast[6]
port 52 nsew signal output
rlabel metal3 s 179200 95208 180000 95328 6 oeast[7]
port 53 nsew signal output
rlabel metal3 s 179200 100648 180000 100768 6 oeast[8]
port 54 nsew signal output
rlabel metal3 s 179200 106088 180000 106208 6 oeast[9]
port 55 nsew signal output
rlabel metal2 s 85486 119200 85542 120000 6 onorth[0]
port 56 nsew signal output
rlabel metal2 s 76562 119200 76618 120000 6 onorth[1]
port 57 nsew signal output
rlabel metal2 s 67638 119200 67694 120000 6 onorth[2]
port 58 nsew signal output
rlabel metal2 s 58714 119200 58770 120000 6 onorth[3]
port 59 nsew signal output
rlabel metal2 s 49790 119200 49846 120000 6 onorth[4]
port 60 nsew signal output
rlabel metal2 s 40866 119200 40922 120000 6 onorth[5]
port 61 nsew signal output
rlabel metal2 s 31942 119200 31998 120000 6 onorth[6]
port 62 nsew signal output
rlabel metal2 s 23018 119200 23074 120000 6 onorth[7]
port 63 nsew signal output
rlabel metal2 s 14094 119200 14150 120000 6 onorth[8]
port 64 nsew signal output
rlabel metal2 s 5170 119200 5226 120000 6 onorth[9]
port 65 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 osouth[0]
port 66 nsew signal output
rlabel metal2 s 110234 0 110290 800 6 osouth[1]
port 67 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 osouth[2]
port 68 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 osouth[3]
port 69 nsew signal output
rlabel metal2 s 134522 0 134578 800 6 osouth[4]
port 70 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 osouth[5]
port 71 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 osouth[6]
port 72 nsew signal output
rlabel metal2 s 158810 0 158866 800 6 osouth[7]
port 73 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 osouth[8]
port 74 nsew signal output
rlabel metal2 s 175002 0 175058 800 6 osouth[9]
port 75 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 owest[0]
port 76 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 owest[1]
port 77 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 owest[2]
port 78 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 owest[3]
port 79 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 owest[4]
port 80 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 owest[5]
port 81 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 owest[6]
port 82 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 owest[7]
port 83 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 owest[8]
port 84 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 owest[9]
port 85 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 reset
port 86 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 87 nsew power bidirectional
rlabel metal5 s 1056 5346 178896 5666 6 vccd1
port 87 nsew power bidirectional
rlabel metal5 s 1056 35982 178896 36302 6 vccd1
port 87 nsew power bidirectional
rlabel metal5 s 1056 66618 178896 66938 6 vccd1
port 87 nsew power bidirectional
rlabel metal5 s 1056 97254 178896 97574 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 88 nsew ground bidirectional
rlabel metal5 s 1056 20664 178896 20984 6 vssd1
port 88 nsew ground bidirectional
rlabel metal5 s 1056 51300 178896 51620 6 vssd1
port 88 nsew ground bidirectional
rlabel metal5 s 1056 81936 178896 82256 6 vssd1
port 88 nsew ground bidirectional
rlabel metal5 s 1056 112572 178896 112892 6 vssd1
port 88 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 36487724
string GDS_FILE /home/alex/chaos_automaton_Summer_2022/openlane/chaos_subarray/runs/22_08_05_16_33/results/signoff/chaos_subarray.magic.gds
string GDS_START 141920
<< end >>

