magic
tech sky130B
magscale 1 2
timestamp 1660324207
<< obsli1 >>
rect 1104 2159 582820 701777
<< obsm1 >>
rect 566 1844 583450 701808
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 572 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 583444 703610
rect 572 536 583444 703464
rect 710 326 1590 536
rect 1814 326 2786 536
rect 3010 326 3982 536
rect 4206 326 5178 536
rect 5402 326 6374 536
rect 6598 326 7570 536
rect 7794 326 8674 536
rect 8898 326 9870 536
rect 10094 326 11066 536
rect 11290 326 12262 536
rect 12486 326 13458 536
rect 13682 326 14654 536
rect 14878 326 15850 536
rect 16074 326 16954 536
rect 17178 326 18150 536
rect 18374 326 19346 536
rect 19570 326 20542 536
rect 20766 326 21738 536
rect 21962 326 22934 536
rect 23158 326 24130 536
rect 24354 326 25234 536
rect 25458 326 26430 536
rect 26654 326 27626 536
rect 27850 326 28822 536
rect 29046 326 30018 536
rect 30242 326 31214 536
rect 31438 326 32318 536
rect 32542 326 33514 536
rect 33738 326 34710 536
rect 34934 326 35906 536
rect 36130 326 37102 536
rect 37326 326 38298 536
rect 38522 326 39494 536
rect 39718 326 40598 536
rect 40822 326 41794 536
rect 42018 326 42990 536
rect 43214 326 44186 536
rect 44410 326 45382 536
rect 45606 326 46578 536
rect 46802 326 47774 536
rect 47998 326 48878 536
rect 49102 326 50074 536
rect 50298 326 51270 536
rect 51494 326 52466 536
rect 52690 326 53662 536
rect 53886 326 54858 536
rect 55082 326 55962 536
rect 56186 326 57158 536
rect 57382 326 58354 536
rect 58578 326 59550 536
rect 59774 326 60746 536
rect 60970 326 61942 536
rect 62166 326 63138 536
rect 63362 326 64242 536
rect 64466 326 65438 536
rect 65662 326 66634 536
rect 66858 326 67830 536
rect 68054 326 69026 536
rect 69250 326 70222 536
rect 70446 326 71418 536
rect 71642 326 72522 536
rect 72746 326 73718 536
rect 73942 326 74914 536
rect 75138 326 76110 536
rect 76334 326 77306 536
rect 77530 326 78502 536
rect 78726 326 79606 536
rect 79830 326 80802 536
rect 81026 326 81998 536
rect 82222 326 83194 536
rect 83418 326 84390 536
rect 84614 326 85586 536
rect 85810 326 86782 536
rect 87006 326 87886 536
rect 88110 326 89082 536
rect 89306 326 90278 536
rect 90502 326 91474 536
rect 91698 326 92670 536
rect 92894 326 93866 536
rect 94090 326 95062 536
rect 95286 326 96166 536
rect 96390 326 97362 536
rect 97586 326 98558 536
rect 98782 326 99754 536
rect 99978 326 100950 536
rect 101174 326 102146 536
rect 102370 326 103250 536
rect 103474 326 104446 536
rect 104670 326 105642 536
rect 105866 326 106838 536
rect 107062 326 108034 536
rect 108258 326 109230 536
rect 109454 326 110426 536
rect 110650 326 111530 536
rect 111754 326 112726 536
rect 112950 326 113922 536
rect 114146 326 115118 536
rect 115342 326 116314 536
rect 116538 326 117510 536
rect 117734 326 118706 536
rect 118930 326 119810 536
rect 120034 326 121006 536
rect 121230 326 122202 536
rect 122426 326 123398 536
rect 123622 326 124594 536
rect 124818 326 125790 536
rect 126014 326 126894 536
rect 127118 326 128090 536
rect 128314 326 129286 536
rect 129510 326 130482 536
rect 130706 326 131678 536
rect 131902 326 132874 536
rect 133098 326 134070 536
rect 134294 326 135174 536
rect 135398 326 136370 536
rect 136594 326 137566 536
rect 137790 326 138762 536
rect 138986 326 139958 536
rect 140182 326 141154 536
rect 141378 326 142350 536
rect 142574 326 143454 536
rect 143678 326 144650 536
rect 144874 326 145846 536
rect 146070 326 147042 536
rect 147266 326 148238 536
rect 148462 326 149434 536
rect 149658 326 150538 536
rect 150762 326 151734 536
rect 151958 326 152930 536
rect 153154 326 154126 536
rect 154350 326 155322 536
rect 155546 326 156518 536
rect 156742 326 157714 536
rect 157938 326 158818 536
rect 159042 326 160014 536
rect 160238 326 161210 536
rect 161434 326 162406 536
rect 162630 326 163602 536
rect 163826 326 164798 536
rect 165022 326 165994 536
rect 166218 326 167098 536
rect 167322 326 168294 536
rect 168518 326 169490 536
rect 169714 326 170686 536
rect 170910 326 171882 536
rect 172106 326 173078 536
rect 173302 326 174182 536
rect 174406 326 175378 536
rect 175602 326 176574 536
rect 176798 326 177770 536
rect 177994 326 178966 536
rect 179190 326 180162 536
rect 180386 326 181358 536
rect 181582 326 182462 536
rect 182686 326 183658 536
rect 183882 326 184854 536
rect 185078 326 186050 536
rect 186274 326 187246 536
rect 187470 326 188442 536
rect 188666 326 189638 536
rect 189862 326 190742 536
rect 190966 326 191938 536
rect 192162 326 193134 536
rect 193358 326 194330 536
rect 194554 326 195526 536
rect 195750 326 196722 536
rect 196946 326 197826 536
rect 198050 326 199022 536
rect 199246 326 200218 536
rect 200442 326 201414 536
rect 201638 326 202610 536
rect 202834 326 203806 536
rect 204030 326 205002 536
rect 205226 326 206106 536
rect 206330 326 207302 536
rect 207526 326 208498 536
rect 208722 326 209694 536
rect 209918 326 210890 536
rect 211114 326 212086 536
rect 212310 326 213282 536
rect 213506 326 214386 536
rect 214610 326 215582 536
rect 215806 326 216778 536
rect 217002 326 217974 536
rect 218198 326 219170 536
rect 219394 326 220366 536
rect 220590 326 221470 536
rect 221694 326 222666 536
rect 222890 326 223862 536
rect 224086 326 225058 536
rect 225282 326 226254 536
rect 226478 326 227450 536
rect 227674 326 228646 536
rect 228870 326 229750 536
rect 229974 326 230946 536
rect 231170 326 232142 536
rect 232366 326 233338 536
rect 233562 326 234534 536
rect 234758 326 235730 536
rect 235954 326 236926 536
rect 237150 326 238030 536
rect 238254 326 239226 536
rect 239450 326 240422 536
rect 240646 326 241618 536
rect 241842 326 242814 536
rect 243038 326 244010 536
rect 244234 326 245114 536
rect 245338 326 246310 536
rect 246534 326 247506 536
rect 247730 326 248702 536
rect 248926 326 249898 536
rect 250122 326 251094 536
rect 251318 326 252290 536
rect 252514 326 253394 536
rect 253618 326 254590 536
rect 254814 326 255786 536
rect 256010 326 256982 536
rect 257206 326 258178 536
rect 258402 326 259374 536
rect 259598 326 260570 536
rect 260794 326 261674 536
rect 261898 326 262870 536
rect 263094 326 264066 536
rect 264290 326 265262 536
rect 265486 326 266458 536
rect 266682 326 267654 536
rect 267878 326 268758 536
rect 268982 326 269954 536
rect 270178 326 271150 536
rect 271374 326 272346 536
rect 272570 326 273542 536
rect 273766 326 274738 536
rect 274962 326 275934 536
rect 276158 326 277038 536
rect 277262 326 278234 536
rect 278458 326 279430 536
rect 279654 326 280626 536
rect 280850 326 281822 536
rect 282046 326 283018 536
rect 283242 326 284214 536
rect 284438 326 285318 536
rect 285542 326 286514 536
rect 286738 326 287710 536
rect 287934 326 288906 536
rect 289130 326 290102 536
rect 290326 326 291298 536
rect 291522 326 292494 536
rect 292718 326 293598 536
rect 293822 326 294794 536
rect 295018 326 295990 536
rect 296214 326 297186 536
rect 297410 326 298382 536
rect 298606 326 299578 536
rect 299802 326 300682 536
rect 300906 326 301878 536
rect 302102 326 303074 536
rect 303298 326 304270 536
rect 304494 326 305466 536
rect 305690 326 306662 536
rect 306886 326 307858 536
rect 308082 326 308962 536
rect 309186 326 310158 536
rect 310382 326 311354 536
rect 311578 326 312550 536
rect 312774 326 313746 536
rect 313970 326 314942 536
rect 315166 326 316138 536
rect 316362 326 317242 536
rect 317466 326 318438 536
rect 318662 326 319634 536
rect 319858 326 320830 536
rect 321054 326 322026 536
rect 322250 326 323222 536
rect 323446 326 324326 536
rect 324550 326 325522 536
rect 325746 326 326718 536
rect 326942 326 327914 536
rect 328138 326 329110 536
rect 329334 326 330306 536
rect 330530 326 331502 536
rect 331726 326 332606 536
rect 332830 326 333802 536
rect 334026 326 334998 536
rect 335222 326 336194 536
rect 336418 326 337390 536
rect 337614 326 338586 536
rect 338810 326 339782 536
rect 340006 326 340886 536
rect 341110 326 342082 536
rect 342306 326 343278 536
rect 343502 326 344474 536
rect 344698 326 345670 536
rect 345894 326 346866 536
rect 347090 326 347970 536
rect 348194 326 349166 536
rect 349390 326 350362 536
rect 350586 326 351558 536
rect 351782 326 352754 536
rect 352978 326 353950 536
rect 354174 326 355146 536
rect 355370 326 356250 536
rect 356474 326 357446 536
rect 357670 326 358642 536
rect 358866 326 359838 536
rect 360062 326 361034 536
rect 361258 326 362230 536
rect 362454 326 363426 536
rect 363650 326 364530 536
rect 364754 326 365726 536
rect 365950 326 366922 536
rect 367146 326 368118 536
rect 368342 326 369314 536
rect 369538 326 370510 536
rect 370734 326 371614 536
rect 371838 326 372810 536
rect 373034 326 374006 536
rect 374230 326 375202 536
rect 375426 326 376398 536
rect 376622 326 377594 536
rect 377818 326 378790 536
rect 379014 326 379894 536
rect 380118 326 381090 536
rect 381314 326 382286 536
rect 382510 326 383482 536
rect 383706 326 384678 536
rect 384902 326 385874 536
rect 386098 326 387070 536
rect 387294 326 388174 536
rect 388398 326 389370 536
rect 389594 326 390566 536
rect 390790 326 391762 536
rect 391986 326 392958 536
rect 393182 326 394154 536
rect 394378 326 395258 536
rect 395482 326 396454 536
rect 396678 326 397650 536
rect 397874 326 398846 536
rect 399070 326 400042 536
rect 400266 326 401238 536
rect 401462 326 402434 536
rect 402658 326 403538 536
rect 403762 326 404734 536
rect 404958 326 405930 536
rect 406154 326 407126 536
rect 407350 326 408322 536
rect 408546 326 409518 536
rect 409742 326 410714 536
rect 410938 326 411818 536
rect 412042 326 413014 536
rect 413238 326 414210 536
rect 414434 326 415406 536
rect 415630 326 416602 536
rect 416826 326 417798 536
rect 418022 326 418902 536
rect 419126 326 420098 536
rect 420322 326 421294 536
rect 421518 326 422490 536
rect 422714 326 423686 536
rect 423910 326 424882 536
rect 425106 326 426078 536
rect 426302 326 427182 536
rect 427406 326 428378 536
rect 428602 326 429574 536
rect 429798 326 430770 536
rect 430994 326 431966 536
rect 432190 326 433162 536
rect 433386 326 434358 536
rect 434582 326 435462 536
rect 435686 326 436658 536
rect 436882 326 437854 536
rect 438078 326 439050 536
rect 439274 326 440246 536
rect 440470 326 441442 536
rect 441666 326 442546 536
rect 442770 326 443742 536
rect 443966 326 444938 536
rect 445162 326 446134 536
rect 446358 326 447330 536
rect 447554 326 448526 536
rect 448750 326 449722 536
rect 449946 326 450826 536
rect 451050 326 452022 536
rect 452246 326 453218 536
rect 453442 326 454414 536
rect 454638 326 455610 536
rect 455834 326 456806 536
rect 457030 326 458002 536
rect 458226 326 459106 536
rect 459330 326 460302 536
rect 460526 326 461498 536
rect 461722 326 462694 536
rect 462918 326 463890 536
rect 464114 326 465086 536
rect 465310 326 466190 536
rect 466414 326 467386 536
rect 467610 326 468582 536
rect 468806 326 469778 536
rect 470002 326 470974 536
rect 471198 326 472170 536
rect 472394 326 473366 536
rect 473590 326 474470 536
rect 474694 326 475666 536
rect 475890 326 476862 536
rect 477086 326 478058 536
rect 478282 326 479254 536
rect 479478 326 480450 536
rect 480674 326 481646 536
rect 481870 326 482750 536
rect 482974 326 483946 536
rect 484170 326 485142 536
rect 485366 326 486338 536
rect 486562 326 487534 536
rect 487758 326 488730 536
rect 488954 326 489834 536
rect 490058 326 491030 536
rect 491254 326 492226 536
rect 492450 326 493422 536
rect 493646 326 494618 536
rect 494842 326 495814 536
rect 496038 326 497010 536
rect 497234 326 498114 536
rect 498338 326 499310 536
rect 499534 326 500506 536
rect 500730 326 501702 536
rect 501926 326 502898 536
rect 503122 326 504094 536
rect 504318 326 505290 536
rect 505514 326 506394 536
rect 506618 326 507590 536
rect 507814 326 508786 536
rect 509010 326 509982 536
rect 510206 326 511178 536
rect 511402 326 512374 536
rect 512598 326 513478 536
rect 513702 326 514674 536
rect 514898 326 515870 536
rect 516094 326 517066 536
rect 517290 326 518262 536
rect 518486 326 519458 536
rect 519682 326 520654 536
rect 520878 326 521758 536
rect 521982 326 522954 536
rect 523178 326 524150 536
rect 524374 326 525346 536
rect 525570 326 526542 536
rect 526766 326 527738 536
rect 527962 326 528934 536
rect 529158 326 530038 536
rect 530262 326 531234 536
rect 531458 326 532430 536
rect 532654 326 533626 536
rect 533850 326 534822 536
rect 535046 326 536018 536
rect 536242 326 537122 536
rect 537346 326 538318 536
rect 538542 326 539514 536
rect 539738 326 540710 536
rect 540934 326 541906 536
rect 542130 326 543102 536
rect 543326 326 544298 536
rect 544522 326 545402 536
rect 545626 326 546598 536
rect 546822 326 547794 536
rect 548018 326 548990 536
rect 549214 326 550186 536
rect 550410 326 551382 536
rect 551606 326 552578 536
rect 552802 326 553682 536
rect 553906 326 554878 536
rect 555102 326 556074 536
rect 556298 326 557270 536
rect 557494 326 558466 536
rect 558690 326 559662 536
rect 559886 326 560766 536
rect 560990 326 561962 536
rect 562186 326 563158 536
rect 563382 326 564354 536
rect 564578 326 565550 536
rect 565774 326 566746 536
rect 566970 326 567942 536
rect 568166 326 569046 536
rect 569270 326 570242 536
rect 570466 326 571438 536
rect 571662 326 572634 536
rect 572858 326 573830 536
rect 574054 326 575026 536
rect 575250 326 576222 536
rect 576446 326 577326 536
rect 577550 326 578522 536
rect 578746 326 579718 536
rect 579942 326 580914 536
rect 581138 326 582110 536
rect 582334 326 583306 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 480 697540 583520 701793
rect 560 697404 583520 697540
rect 560 697140 583440 697404
rect 480 697004 583440 697140
rect 480 684484 583520 697004
rect 560 684084 583520 684484
rect 480 684076 583520 684084
rect 480 683676 583440 684076
rect 480 671428 583520 683676
rect 560 671028 583520 671428
rect 480 670884 583520 671028
rect 480 670484 583440 670884
rect 480 658372 583520 670484
rect 560 657972 583520 658372
rect 480 657556 583520 657972
rect 480 657156 583440 657556
rect 480 645316 583520 657156
rect 560 644916 583520 645316
rect 480 644228 583520 644916
rect 480 643828 583440 644228
rect 480 632260 583520 643828
rect 560 631860 583520 632260
rect 480 631036 583520 631860
rect 480 630636 583440 631036
rect 480 619340 583520 630636
rect 560 618940 583520 619340
rect 480 617708 583520 618940
rect 480 617308 583440 617708
rect 480 606284 583520 617308
rect 560 605884 583520 606284
rect 480 604380 583520 605884
rect 480 603980 583440 604380
rect 480 593228 583520 603980
rect 560 592828 583520 593228
rect 480 591188 583520 592828
rect 480 590788 583440 591188
rect 480 580172 583520 590788
rect 560 579772 583520 580172
rect 480 577860 583520 579772
rect 480 577460 583440 577860
rect 480 567116 583520 577460
rect 560 566716 583520 567116
rect 480 564532 583520 566716
rect 480 564132 583440 564532
rect 480 554060 583520 564132
rect 560 553660 583520 554060
rect 480 551340 583520 553660
rect 480 550940 583440 551340
rect 480 541004 583520 550940
rect 560 540604 583520 541004
rect 480 538012 583520 540604
rect 480 537612 583440 538012
rect 480 528084 583520 537612
rect 560 527684 583520 528084
rect 480 524684 583520 527684
rect 480 524284 583440 524684
rect 480 515028 583520 524284
rect 560 514628 583520 515028
rect 480 511492 583520 514628
rect 480 511092 583440 511492
rect 480 501972 583520 511092
rect 560 501572 583520 501972
rect 480 498164 583520 501572
rect 480 497764 583440 498164
rect 480 488916 583520 497764
rect 560 488516 583520 488916
rect 480 484836 583520 488516
rect 480 484436 583440 484836
rect 480 475860 583520 484436
rect 560 475460 583520 475860
rect 480 471644 583520 475460
rect 480 471244 583440 471644
rect 480 462804 583520 471244
rect 560 462404 583520 462804
rect 480 458316 583520 462404
rect 480 457916 583440 458316
rect 480 449748 583520 457916
rect 560 449348 583520 449748
rect 480 444988 583520 449348
rect 480 444588 583440 444988
rect 480 436828 583520 444588
rect 560 436428 583520 436828
rect 480 431796 583520 436428
rect 480 431396 583440 431796
rect 480 423772 583520 431396
rect 560 423372 583520 423772
rect 480 418468 583520 423372
rect 480 418068 583440 418468
rect 480 410716 583520 418068
rect 560 410316 583520 410716
rect 480 405140 583520 410316
rect 480 404740 583440 405140
rect 480 397660 583520 404740
rect 560 397260 583520 397660
rect 480 391948 583520 397260
rect 480 391548 583440 391948
rect 480 384604 583520 391548
rect 560 384204 583520 384604
rect 480 378620 583520 384204
rect 480 378220 583440 378620
rect 480 371548 583520 378220
rect 560 371148 583520 371548
rect 480 365292 583520 371148
rect 480 364892 583440 365292
rect 480 358628 583520 364892
rect 560 358228 583520 358628
rect 480 352100 583520 358228
rect 480 351700 583440 352100
rect 480 345572 583520 351700
rect 560 345172 583520 345572
rect 480 338772 583520 345172
rect 480 338372 583440 338772
rect 480 332516 583520 338372
rect 560 332116 583520 332516
rect 480 325444 583520 332116
rect 480 325044 583440 325444
rect 480 319460 583520 325044
rect 560 319060 583520 319460
rect 480 312252 583520 319060
rect 480 311852 583440 312252
rect 480 306404 583520 311852
rect 560 306004 583520 306404
rect 480 298924 583520 306004
rect 480 298524 583440 298924
rect 480 293348 583520 298524
rect 560 292948 583520 293348
rect 480 285596 583520 292948
rect 480 285196 583440 285596
rect 480 280292 583520 285196
rect 560 279892 583520 280292
rect 480 272404 583520 279892
rect 480 272004 583440 272404
rect 480 267372 583520 272004
rect 560 266972 583520 267372
rect 480 259076 583520 266972
rect 480 258676 583440 259076
rect 480 254316 583520 258676
rect 560 253916 583520 254316
rect 480 245748 583520 253916
rect 480 245348 583440 245748
rect 480 241260 583520 245348
rect 560 240860 583520 241260
rect 480 232556 583520 240860
rect 480 232156 583440 232556
rect 480 228204 583520 232156
rect 560 227804 583520 228204
rect 480 219228 583520 227804
rect 480 218828 583440 219228
rect 480 215148 583520 218828
rect 560 214748 583520 215148
rect 480 205900 583520 214748
rect 480 205500 583440 205900
rect 480 202092 583520 205500
rect 560 201692 583520 202092
rect 480 192708 583520 201692
rect 480 192308 583440 192708
rect 480 189036 583520 192308
rect 560 188636 583520 189036
rect 480 179380 583520 188636
rect 480 178980 583440 179380
rect 480 176116 583520 178980
rect 560 175716 583520 176116
rect 480 166052 583520 175716
rect 480 165652 583440 166052
rect 480 163060 583520 165652
rect 560 162660 583520 163060
rect 480 152860 583520 162660
rect 480 152460 583440 152860
rect 480 150004 583520 152460
rect 560 149604 583520 150004
rect 480 139532 583520 149604
rect 480 139132 583440 139532
rect 480 136948 583520 139132
rect 560 136548 583520 136948
rect 480 126204 583520 136548
rect 480 125804 583440 126204
rect 480 123892 583520 125804
rect 560 123492 583520 123892
rect 480 113012 583520 123492
rect 480 112612 583440 113012
rect 480 110836 583520 112612
rect 560 110436 583520 110836
rect 480 99684 583520 110436
rect 480 99284 583440 99684
rect 480 97780 583520 99284
rect 560 97380 583520 97780
rect 480 86356 583520 97380
rect 480 85956 583440 86356
rect 480 84860 583520 85956
rect 560 84460 583520 84860
rect 480 73164 583520 84460
rect 480 72764 583440 73164
rect 480 71804 583520 72764
rect 560 71404 583520 71804
rect 480 59836 583520 71404
rect 480 59436 583440 59836
rect 480 58748 583520 59436
rect 560 58348 583520 58748
rect 480 46508 583520 58348
rect 480 46108 583440 46508
rect 480 45692 583520 46108
rect 560 45292 583520 45692
rect 480 33316 583520 45292
rect 480 32916 583440 33316
rect 480 32636 583520 32916
rect 560 32236 583520 32636
rect 480 19988 583520 32236
rect 480 19588 583440 19988
rect 480 19580 583520 19588
rect 560 19180 583520 19580
rect 480 6796 583520 19180
rect 480 6660 583440 6796
rect 560 6396 583440 6660
rect 560 6260 583520 6396
rect 480 2143 583520 6260
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 4058 -7654 4678 711590
rect 7898 -7654 8518 711590
rect 34778 687000 35398 711590
rect 38618 687000 39238 711590
rect 65498 687000 66118 711590
rect 69338 687000 69958 711590
rect 96218 687000 96838 711590
rect 100058 687000 100678 711590
rect 126938 687000 127558 711590
rect 130778 687000 131398 711590
rect 157658 687000 158278 711590
rect 161498 687000 162118 711590
rect 188378 687000 188998 711590
rect 34778 550000 35398 566000
rect 38618 550000 39238 566000
rect 65498 550000 66118 566000
rect 69338 550000 69958 566000
rect 96218 550000 96838 566000
rect 100058 550000 100678 566000
rect 126938 550000 127558 566000
rect 130778 550000 131398 566000
rect 157658 550000 158278 566000
rect 161498 550000 162118 566000
rect 188378 550000 188998 566000
rect 34778 413000 35398 429000
rect 38618 413000 39238 429000
rect 65498 413000 66118 429000
rect 69338 413000 69958 429000
rect 96218 413000 96838 429000
rect 100058 413000 100678 429000
rect 126938 413000 127558 429000
rect 130778 413000 131398 429000
rect 157658 413000 158278 429000
rect 161498 413000 162118 429000
rect 188378 413000 188998 429000
rect 34778 276000 35398 292000
rect 38618 276000 39238 292000
rect 65498 276000 66118 292000
rect 69338 276000 69958 292000
rect 96218 276000 96838 292000
rect 100058 276000 100678 292000
rect 126938 276000 127558 292000
rect 130778 276000 131398 292000
rect 157658 276000 158278 292000
rect 161498 276000 162118 292000
rect 188378 276000 188998 292000
rect 34778 139000 35398 155000
rect 38618 139000 39238 155000
rect 65498 139000 66118 155000
rect 69338 139000 69958 155000
rect 96218 139000 96838 155000
rect 100058 139000 100678 155000
rect 126938 139000 127558 155000
rect 130778 139000 131398 155000
rect 157658 139000 158278 155000
rect 161498 139000 162118 155000
rect 188378 139000 188998 155000
rect 34778 -7654 35398 18000
rect 38618 -7654 39238 18000
rect 65498 -7654 66118 18000
rect 69338 -7654 69958 18000
rect 96218 -7654 96838 18000
rect 100058 -7654 100678 18000
rect 126938 -7654 127558 18000
rect 130778 -7654 131398 18000
rect 157658 -7654 158278 18000
rect 161498 -7654 162118 18000
rect 188378 -7654 188998 18000
rect 192218 -7654 192838 711590
rect 198134 565712 198754 687664
rect 219098 687000 219718 711590
rect 222938 687000 223558 711590
rect 249818 687000 250438 711590
rect 253658 687000 254278 711590
rect 280538 687000 281158 711590
rect 284378 687000 284998 711590
rect 311258 687000 311878 711590
rect 315098 687000 315718 711590
rect 341978 687000 342598 711590
rect 345818 687000 346438 711590
rect 372698 687000 373318 711590
rect 198134 428624 198754 550576
rect 219098 550000 219718 566000
rect 222938 550000 223558 566000
rect 249818 550000 250438 566000
rect 253658 550000 254278 566000
rect 280538 550000 281158 566000
rect 284378 550000 284998 566000
rect 311258 550000 311878 566000
rect 315098 550000 315718 566000
rect 341978 550000 342598 566000
rect 345818 550000 346438 566000
rect 372698 550000 373318 566000
rect 198134 291536 198754 413488
rect 219098 413000 219718 429000
rect 222938 413000 223558 429000
rect 249818 413000 250438 429000
rect 253658 413000 254278 429000
rect 280538 413000 281158 429000
rect 284378 413000 284998 429000
rect 311258 413000 311878 429000
rect 315098 413000 315718 429000
rect 341978 413000 342598 429000
rect 345818 413000 346438 429000
rect 372698 413000 373318 429000
rect 198134 154448 198754 276400
rect 219098 276000 219718 292000
rect 222938 276000 223558 292000
rect 249818 276000 250438 292000
rect 253658 276000 254278 292000
rect 280538 276000 281158 292000
rect 284378 276000 284998 292000
rect 311258 276000 311878 292000
rect 315098 276000 315718 292000
rect 341978 276000 342598 292000
rect 345818 276000 346438 292000
rect 372698 276000 373318 292000
rect 198134 17360 198754 139312
rect 219098 139000 219718 155000
rect 222938 139000 223558 155000
rect 249818 139000 250438 155000
rect 253658 139000 254278 155000
rect 280538 139000 281158 155000
rect 284378 139000 284998 155000
rect 311258 139000 311878 155000
rect 315098 139000 315718 155000
rect 341978 139000 342598 155000
rect 345818 139000 346438 155000
rect 372698 139000 373318 155000
rect 219098 -7654 219718 18000
rect 222938 -7654 223558 18000
rect 249818 -7654 250438 18000
rect 253658 -7654 254278 18000
rect 280538 -7654 281158 18000
rect 284378 -7654 284998 18000
rect 311258 -7654 311878 18000
rect 315098 -7654 315718 18000
rect 341978 -7654 342598 18000
rect 345818 -7654 346438 18000
rect 372698 -7654 373318 18000
rect 376538 -7654 377158 711590
rect 385262 565712 385882 687664
rect 403418 687000 404038 711590
rect 407258 687000 407878 711590
rect 434138 687000 434758 711590
rect 437978 687000 438598 711590
rect 464858 687000 465478 711590
rect 468698 687000 469318 711590
rect 495578 687000 496198 711590
rect 499418 687000 500038 711590
rect 526298 687000 526918 711590
rect 530138 687000 530758 711590
rect 557018 687000 557638 711590
rect 560858 687000 561478 711590
rect 385262 428624 385882 550576
rect 403418 550000 404038 566000
rect 407258 550000 407878 566000
rect 434138 550000 434758 566000
rect 437978 550000 438598 566000
rect 464858 550000 465478 566000
rect 468698 550000 469318 566000
rect 495578 550000 496198 566000
rect 499418 550000 500038 566000
rect 526298 550000 526918 566000
rect 530138 550000 530758 566000
rect 557018 550000 557638 566000
rect 560858 550000 561478 566000
rect 571102 565168 571722 687664
rect 574966 565168 575586 687664
rect 385262 291536 385882 413488
rect 403418 413000 404038 429000
rect 407258 413000 407878 429000
rect 434138 413000 434758 429000
rect 437978 413000 438598 429000
rect 464858 413000 465478 429000
rect 468698 413000 469318 429000
rect 495578 413000 496198 429000
rect 499418 413000 500038 429000
rect 526298 413000 526918 429000
rect 530138 413000 530758 429000
rect 557018 413000 557638 429000
rect 560858 413000 561478 429000
rect 571102 428080 571722 551120
rect 574966 428080 575586 551120
rect 385262 154448 385882 276400
rect 403418 276000 404038 292000
rect 407258 276000 407878 292000
rect 434138 276000 434758 292000
rect 437978 276000 438598 292000
rect 464858 276000 465478 292000
rect 468698 276000 469318 292000
rect 495578 276000 496198 292000
rect 499418 276000 500038 292000
rect 526298 276000 526918 292000
rect 530138 276000 530758 292000
rect 557018 276000 557638 292000
rect 560858 276000 561478 292000
rect 571102 290992 571722 414032
rect 574966 290992 575586 414032
rect 385262 17360 385882 139312
rect 403418 139000 404038 155000
rect 407258 139000 407878 155000
rect 434138 139000 434758 155000
rect 437978 139000 438598 155000
rect 464858 139000 465478 155000
rect 468698 139000 469318 155000
rect 495578 139000 496198 155000
rect 499418 139000 500038 155000
rect 526298 139000 526918 155000
rect 530138 139000 530758 155000
rect 557018 139000 557638 155000
rect 560858 139000 561478 155000
rect 571102 153904 571722 276944
rect 574966 153904 575586 276944
rect 403418 -7654 404038 18000
rect 407258 -7654 407878 18000
rect 434138 -7654 434758 18000
rect 437978 -7654 438598 18000
rect 464858 -7654 465478 18000
rect 468698 -7654 469318 18000
rect 495578 -7654 496198 18000
rect 499418 -7654 500038 18000
rect 526298 -7654 526918 18000
rect 530138 -7654 530758 18000
rect 557018 -7654 557638 18000
rect 560858 -7654 561478 18000
rect 571102 17360 571722 139856
rect 574966 17360 575586 139856
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 2366 2347 3978 688533
rect 4758 2347 7818 688533
rect 8598 686920 34698 688533
rect 35478 686920 38538 688533
rect 39318 686920 65418 688533
rect 66198 686920 69258 688533
rect 70038 686920 96138 688533
rect 96918 686920 99978 688533
rect 100758 686920 126858 688533
rect 127638 686920 130698 688533
rect 131478 686920 157578 688533
rect 158358 686920 161418 688533
rect 162198 686920 188298 688533
rect 189078 686920 192138 688533
rect 8598 566080 192138 686920
rect 8598 549920 34698 566080
rect 35478 549920 38538 566080
rect 39318 549920 65418 566080
rect 66198 549920 69258 566080
rect 70038 549920 96138 566080
rect 96918 549920 99978 566080
rect 100758 549920 126858 566080
rect 127638 549920 130698 566080
rect 131478 549920 157578 566080
rect 158358 549920 161418 566080
rect 162198 549920 188298 566080
rect 189078 549920 192138 566080
rect 8598 429080 192138 549920
rect 8598 412920 34698 429080
rect 35478 412920 38538 429080
rect 39318 412920 65418 429080
rect 66198 412920 69258 429080
rect 70038 412920 96138 429080
rect 96918 412920 99978 429080
rect 100758 412920 126858 429080
rect 127638 412920 130698 429080
rect 131478 412920 157578 429080
rect 158358 412920 161418 429080
rect 162198 412920 188298 429080
rect 189078 412920 192138 429080
rect 8598 292080 192138 412920
rect 8598 275920 34698 292080
rect 35478 275920 38538 292080
rect 39318 275920 65418 292080
rect 66198 275920 69258 292080
rect 70038 275920 96138 292080
rect 96918 275920 99978 292080
rect 100758 275920 126858 292080
rect 127638 275920 130698 292080
rect 131478 275920 157578 292080
rect 158358 275920 161418 292080
rect 162198 275920 188298 292080
rect 189078 275920 192138 292080
rect 8598 155080 192138 275920
rect 8598 138920 34698 155080
rect 35478 138920 38538 155080
rect 39318 138920 65418 155080
rect 66198 138920 69258 155080
rect 70038 138920 96138 155080
rect 96918 138920 99978 155080
rect 100758 138920 126858 155080
rect 127638 138920 130698 155080
rect 131478 138920 157578 155080
rect 158358 138920 161418 155080
rect 162198 138920 188298 155080
rect 189078 138920 192138 155080
rect 8598 18080 192138 138920
rect 8598 2347 34698 18080
rect 35478 2347 38538 18080
rect 39318 2347 65418 18080
rect 66198 2347 69258 18080
rect 70038 2347 96138 18080
rect 96918 2347 99978 18080
rect 100758 2347 126858 18080
rect 127638 2347 130698 18080
rect 131478 2347 157578 18080
rect 158358 2347 161418 18080
rect 162198 2347 188298 18080
rect 189078 2347 192138 18080
rect 192918 687744 219018 688533
rect 192918 565632 198054 687744
rect 198834 686920 219018 687744
rect 219798 686920 222858 688533
rect 223638 686920 249738 688533
rect 250518 686920 253578 688533
rect 254358 686920 280458 688533
rect 281238 686920 284298 688533
rect 285078 686920 311178 688533
rect 311958 686920 315018 688533
rect 315798 686920 341898 688533
rect 342678 686920 345738 688533
rect 346518 686920 372618 688533
rect 373398 686920 376458 688533
rect 198834 566080 376458 686920
rect 198834 565632 219018 566080
rect 192918 550656 219018 565632
rect 192918 428544 198054 550656
rect 198834 549920 219018 550656
rect 219798 549920 222858 566080
rect 223638 549920 249738 566080
rect 250518 549920 253578 566080
rect 254358 549920 280458 566080
rect 281238 549920 284298 566080
rect 285078 549920 311178 566080
rect 311958 549920 315018 566080
rect 315798 549920 341898 566080
rect 342678 549920 345738 566080
rect 346518 549920 372618 566080
rect 373398 549920 376458 566080
rect 198834 429080 376458 549920
rect 198834 428544 219018 429080
rect 192918 413568 219018 428544
rect 192918 291456 198054 413568
rect 198834 412920 219018 413568
rect 219798 412920 222858 429080
rect 223638 412920 249738 429080
rect 250518 412920 253578 429080
rect 254358 412920 280458 429080
rect 281238 412920 284298 429080
rect 285078 412920 311178 429080
rect 311958 412920 315018 429080
rect 315798 412920 341898 429080
rect 342678 412920 345738 429080
rect 346518 412920 372618 429080
rect 373398 412920 376458 429080
rect 198834 292080 376458 412920
rect 198834 291456 219018 292080
rect 192918 276480 219018 291456
rect 192918 154368 198054 276480
rect 198834 275920 219018 276480
rect 219798 275920 222858 292080
rect 223638 275920 249738 292080
rect 250518 275920 253578 292080
rect 254358 275920 280458 292080
rect 281238 275920 284298 292080
rect 285078 275920 311178 292080
rect 311958 275920 315018 292080
rect 315798 275920 341898 292080
rect 342678 275920 345738 292080
rect 346518 275920 372618 292080
rect 373398 275920 376458 292080
rect 198834 155080 376458 275920
rect 198834 154368 219018 155080
rect 192918 139392 219018 154368
rect 192918 17280 198054 139392
rect 198834 138920 219018 139392
rect 219798 138920 222858 155080
rect 223638 138920 249738 155080
rect 250518 138920 253578 155080
rect 254358 138920 280458 155080
rect 281238 138920 284298 155080
rect 285078 138920 311178 155080
rect 311958 138920 315018 155080
rect 315798 138920 341898 155080
rect 342678 138920 345738 155080
rect 346518 138920 372618 155080
rect 373398 138920 376458 155080
rect 198834 18080 376458 138920
rect 198834 17280 219018 18080
rect 192918 2347 219018 17280
rect 219798 2347 222858 18080
rect 223638 2347 249738 18080
rect 250518 2347 253578 18080
rect 254358 2347 280458 18080
rect 281238 2347 284298 18080
rect 285078 2347 311178 18080
rect 311958 2347 315018 18080
rect 315798 2347 341898 18080
rect 342678 2347 345738 18080
rect 346518 2347 372618 18080
rect 373398 2347 376458 18080
rect 377238 687744 403338 688533
rect 377238 565632 385182 687744
rect 385962 686920 403338 687744
rect 404118 686920 407178 688533
rect 407958 686920 434058 688533
rect 434838 686920 437898 688533
rect 438678 686920 464778 688533
rect 465558 686920 468618 688533
rect 469398 686920 495498 688533
rect 496278 686920 499338 688533
rect 500118 686920 526218 688533
rect 526998 686920 530058 688533
rect 530838 686920 556938 688533
rect 557718 686920 560778 688533
rect 561558 687744 581098 688533
rect 561558 686920 571022 687744
rect 385962 566080 571022 686920
rect 385962 565632 403338 566080
rect 377238 550656 403338 565632
rect 377238 428544 385182 550656
rect 385962 549920 403338 550656
rect 404118 549920 407178 566080
rect 407958 549920 434058 566080
rect 434838 549920 437898 566080
rect 438678 549920 464778 566080
rect 465558 549920 468618 566080
rect 469398 549920 495498 566080
rect 496278 549920 499338 566080
rect 500118 549920 526218 566080
rect 526998 549920 530058 566080
rect 530838 549920 556938 566080
rect 557718 549920 560778 566080
rect 561558 565088 571022 566080
rect 571802 565088 574886 687744
rect 575666 565088 581098 687744
rect 561558 551200 581098 565088
rect 561558 549920 571022 551200
rect 385962 429080 571022 549920
rect 385962 428544 403338 429080
rect 377238 413568 403338 428544
rect 377238 291456 385182 413568
rect 385962 412920 403338 413568
rect 404118 412920 407178 429080
rect 407958 412920 434058 429080
rect 434838 412920 437898 429080
rect 438678 412920 464778 429080
rect 465558 412920 468618 429080
rect 469398 412920 495498 429080
rect 496278 412920 499338 429080
rect 500118 412920 526218 429080
rect 526998 412920 530058 429080
rect 530838 412920 556938 429080
rect 557718 412920 560778 429080
rect 561558 428000 571022 429080
rect 571802 428000 574886 551200
rect 575666 428000 581098 551200
rect 561558 414112 581098 428000
rect 561558 412920 571022 414112
rect 385962 292080 571022 412920
rect 385962 291456 403338 292080
rect 377238 276480 403338 291456
rect 377238 154368 385182 276480
rect 385962 275920 403338 276480
rect 404118 275920 407178 292080
rect 407958 275920 434058 292080
rect 434838 275920 437898 292080
rect 438678 275920 464778 292080
rect 465558 275920 468618 292080
rect 469398 275920 495498 292080
rect 496278 275920 499338 292080
rect 500118 275920 526218 292080
rect 526998 275920 530058 292080
rect 530838 275920 556938 292080
rect 557718 275920 560778 292080
rect 561558 290912 571022 292080
rect 571802 290912 574886 414112
rect 575666 290912 581098 414112
rect 561558 277024 581098 290912
rect 561558 275920 571022 277024
rect 385962 155080 571022 275920
rect 385962 154368 403338 155080
rect 377238 139392 403338 154368
rect 377238 17280 385182 139392
rect 385962 138920 403338 139392
rect 404118 138920 407178 155080
rect 407958 138920 434058 155080
rect 434838 138920 437898 155080
rect 438678 138920 464778 155080
rect 465558 138920 468618 155080
rect 469398 138920 495498 155080
rect 496278 138920 499338 155080
rect 500118 138920 526218 155080
rect 526998 138920 530058 155080
rect 530838 138920 556938 155080
rect 557718 138920 560778 155080
rect 561558 153824 571022 155080
rect 571802 153824 574886 277024
rect 575666 153824 581098 277024
rect 561558 139936 581098 153824
rect 561558 138920 571022 139936
rect 385962 18080 571022 138920
rect 385962 17280 403338 18080
rect 377238 2347 403338 17280
rect 404118 2347 407178 18080
rect 407958 2347 434058 18080
rect 434838 2347 437898 18080
rect 438678 2347 464778 18080
rect 465558 2347 468618 18080
rect 469398 2347 495498 18080
rect 496278 2347 499338 18080
rect 500118 2347 526218 18080
rect 526998 2347 530058 18080
rect 530838 2347 556938 18080
rect 557718 2347 560778 18080
rect 561558 17280 571022 18080
rect 571802 17280 574886 139936
rect 575666 17280 581098 139936
rect 561558 2347 581098 17280
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 683017 592650 683637
rect -8726 679188 592650 679808
rect -8726 652381 592650 653001
rect -8726 648552 592650 649172
rect -8726 621745 592650 622365
rect -8726 617916 592650 618536
rect -8726 591109 592650 591729
rect -8726 587280 592650 587900
rect -8726 560473 592650 561093
rect -8726 556644 592650 557264
rect -8726 529837 592650 530457
rect -8726 526008 592650 526628
rect -8726 499201 592650 499821
rect -8726 495372 592650 495992
rect -8726 468565 592650 469185
rect -8726 464736 592650 465356
rect -8726 437929 592650 438549
rect -8726 434100 592650 434720
rect 4058 422990 582868 423610
rect 4058 418910 582868 419530
rect -8726 407293 592650 407913
rect -8726 403464 592650 404084
rect -8726 376657 592650 377277
rect -8726 372828 592650 373448
rect -8726 346021 592650 346641
rect -8726 342192 592650 342812
rect -8726 315385 592650 316005
rect -8726 311556 592650 312176
rect -8726 284749 592650 285369
rect -8726 280920 592650 281540
rect -8726 254113 592650 254733
rect -8726 250284 592650 250904
rect -8726 223477 592650 224097
rect -8726 219648 592650 220268
rect -8726 192841 592650 193461
rect -8726 189012 592650 189632
rect -8726 162205 592650 162825
rect -8726 158376 592650 158996
rect 4058 148950 582868 149570
rect 4058 144870 582868 145490
rect -8726 131569 592650 132189
rect -8726 127740 592650 128360
rect -8726 100933 592650 101553
rect -8726 97104 592650 97724
rect -8726 70297 592650 70917
rect -8726 66468 592650 67088
rect -8726 39661 592650 40281
rect -8726 35832 592650 36452
rect -8726 9025 592650 9645
rect -8726 5196 592650 5816
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< obsm5 >>
rect 2324 618856 581140 619300
rect 2324 592049 581140 617596
rect 2324 588220 581140 590789
rect 2324 561413 581140 586960
rect 2324 557584 581140 560153
rect 2324 530777 581140 556324
rect 2324 526948 581140 529517
rect 2324 500141 581140 525688
rect 2324 496312 581140 498881
rect 2324 469505 581140 495052
rect 2324 465676 581140 468245
rect 2324 438869 581140 464416
rect 2324 435040 581140 437609
rect 2324 423930 581140 433780
rect 2324 422670 3738 423930
rect 2324 419850 581140 422670
rect 2324 418590 3738 419850
rect 2324 408233 581140 418590
rect 2324 404404 581140 406973
rect 2324 377597 581140 403144
rect 2324 373768 581140 376337
rect 2324 346961 581140 372508
rect 2324 343132 581140 345701
rect 2324 316325 581140 341872
rect 2324 312496 581140 315065
rect 2324 285689 581140 311236
rect 2324 281860 581140 284429
rect 2324 255053 581140 280600
rect 2324 251224 581140 253793
rect 2324 224417 581140 249964
rect 2324 220588 581140 223157
rect 2324 193781 581140 219328
rect 2324 189952 581140 192521
rect 2324 163145 581140 188692
rect 2324 159316 581140 161885
rect 2324 149890 581140 158056
rect 2324 148630 3738 149890
rect 2324 145810 581140 148630
rect 2324 144550 3738 145810
rect 2324 132509 581140 144550
rect 2324 128680 581140 131249
rect 2324 101873 581140 127420
rect 2324 98044 581140 100613
rect 2324 71237 581140 96784
rect 2324 67408 581140 69977
rect 2324 40601 581140 66148
rect 2324 36772 581140 39341
rect 2324 9965 581140 35512
rect 2324 6136 581140 8705
rect 2324 3580 581140 4876
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 7898 -7654 8518 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 38618 -7654 39238 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 38618 139000 39238 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 38618 276000 39238 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 38618 413000 39238 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 38618 550000 39238 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 38618 687000 39238 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 69338 -7654 69958 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 69338 139000 69958 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 69338 276000 69958 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 69338 413000 69958 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 69338 550000 69958 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 69338 687000 69958 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 100058 -7654 100678 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 100058 139000 100678 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 100058 276000 100678 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 100058 413000 100678 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 100058 550000 100678 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 100058 687000 100678 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 130778 -7654 131398 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 130778 139000 131398 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 130778 276000 131398 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 130778 413000 131398 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 130778 550000 131398 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 130778 687000 131398 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 161498 -7654 162118 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 161498 139000 162118 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 161498 276000 162118 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 161498 413000 162118 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 161498 550000 162118 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 161498 687000 162118 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 192218 -7654 192838 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 222938 -7654 223558 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 222938 139000 223558 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 222938 276000 223558 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 222938 413000 223558 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 222938 550000 223558 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 222938 687000 223558 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253658 -7654 254278 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253658 139000 254278 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253658 276000 254278 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253658 413000 254278 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253658 550000 254278 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253658 687000 254278 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 284378 -7654 284998 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 284378 139000 284998 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 284378 276000 284998 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 284378 413000 284998 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 284378 550000 284998 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 284378 687000 284998 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 315098 -7654 315718 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 315098 139000 315718 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 315098 276000 315718 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 315098 413000 315718 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 315098 550000 315718 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 315098 687000 315718 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 345818 -7654 346438 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 345818 139000 346438 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 345818 276000 346438 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 345818 413000 346438 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 345818 550000 346438 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 345818 687000 346438 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 376538 -7654 377158 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 407258 -7654 407878 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 407258 139000 407878 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 407258 276000 407878 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 407258 413000 407878 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 407258 550000 407878 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 407258 687000 407878 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 437978 -7654 438598 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 437978 139000 438598 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 437978 276000 438598 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 437978 413000 438598 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 437978 550000 438598 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 437978 687000 438598 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 468698 -7654 469318 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 468698 139000 469318 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 468698 276000 469318 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 468698 413000 469318 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 468698 550000 469318 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 468698 687000 469318 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 499418 -7654 500038 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 499418 139000 500038 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 499418 276000 500038 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 499418 413000 500038 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 499418 550000 500038 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 499418 687000 500038 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 530138 -7654 530758 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 530138 139000 530758 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 530138 276000 530758 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 530138 413000 530758 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 530138 550000 530758 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 530138 687000 530758 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 560858 -7654 561478 18000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 560858 139000 561478 155000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 560858 276000 561478 292000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 560858 413000 561478 429000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 560858 550000 561478 566000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 560858 687000 561478 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 9025 592650 9645 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 39661 592650 40281 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 70297 592650 70917 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 100933 592650 101553 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 131569 592650 132189 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 162205 592650 162825 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 192841 592650 193461 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 223477 592650 224097 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 254113 592650 254733 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 284749 592650 285369 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 315385 592650 316005 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 346021 592650 346641 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 376657 592650 377277 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 407293 592650 407913 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 437929 592650 438549 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 468565 592650 469185 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 499201 592650 499821 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 529837 592650 530457 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 560473 592650 561093 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 591109 592650 591729 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 621745 592650 622365 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 652381 592650 653001 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 683017 592650 683637 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 571102 290992 571722 414032 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 571102 428080 571722 551120 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 571102 17360 571722 139856 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 571102 153904 571722 276944 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 571102 565168 571722 687664 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 4058 144870 582868 145490 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 4058 418910 582868 419530 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 4058 -7654 4678 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 34778 -7654 35398 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 34778 139000 35398 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 34778 276000 35398 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 34778 413000 35398 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 34778 550000 35398 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 34778 687000 35398 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65498 -7654 66118 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65498 139000 66118 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65498 276000 66118 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65498 413000 66118 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65498 550000 66118 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65498 687000 66118 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 96218 -7654 96838 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 96218 139000 96838 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 96218 276000 96838 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 96218 413000 96838 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 96218 550000 96838 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 96218 687000 96838 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126938 -7654 127558 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126938 139000 127558 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126938 276000 127558 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126938 413000 127558 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126938 550000 127558 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126938 687000 127558 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 157658 -7654 158278 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 157658 139000 158278 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 157658 276000 158278 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 157658 413000 158278 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 157658 550000 158278 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 157658 687000 158278 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188378 -7654 188998 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188378 139000 188998 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188378 276000 188998 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188378 413000 188998 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188378 550000 188998 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188378 687000 188998 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 219098 -7654 219718 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 219098 139000 219718 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 219098 276000 219718 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 219098 413000 219718 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 219098 550000 219718 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 219098 687000 219718 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 249818 -7654 250438 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 249818 139000 250438 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 249818 276000 250438 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 249818 413000 250438 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 249818 550000 250438 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 249818 687000 250438 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 280538 -7654 281158 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 280538 139000 281158 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 280538 276000 281158 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 280538 413000 281158 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 280538 550000 281158 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 280538 687000 281158 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 311258 -7654 311878 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 311258 139000 311878 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 311258 276000 311878 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 311258 413000 311878 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 311258 550000 311878 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 311258 687000 311878 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 341978 -7654 342598 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 341978 139000 342598 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 341978 276000 342598 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 341978 413000 342598 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 341978 550000 342598 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 341978 687000 342598 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 372698 -7654 373318 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 372698 139000 373318 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 372698 276000 373318 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 372698 413000 373318 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 372698 550000 373318 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 372698 687000 373318 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 403418 -7654 404038 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 403418 139000 404038 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 403418 276000 404038 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 403418 413000 404038 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 403418 550000 404038 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 403418 687000 404038 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 434138 -7654 434758 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 434138 139000 434758 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 434138 276000 434758 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 434138 413000 434758 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 434138 550000 434758 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 434138 687000 434758 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 464858 -7654 465478 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 464858 139000 465478 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 464858 276000 465478 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 464858 413000 465478 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 464858 550000 465478 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 464858 687000 465478 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 495578 -7654 496198 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 495578 139000 496198 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 495578 276000 496198 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 495578 413000 496198 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 495578 550000 496198 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 495578 687000 496198 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 526298 -7654 526918 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 526298 139000 526918 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 526298 276000 526918 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 526298 413000 526918 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 526298 550000 526918 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 526298 687000 526918 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 557018 -7654 557638 18000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 557018 139000 557638 155000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 557018 276000 557638 292000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 557018 413000 557638 429000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 557018 550000 557638 566000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 557018 687000 557638 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 5196 592650 5816 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 35832 592650 36452 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 66468 592650 67088 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 97104 592650 97724 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 127740 592650 128360 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 158376 592650 158996 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 189012 592650 189632 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 219648 592650 220268 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 250284 592650 250904 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 280920 592650 281540 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 311556 592650 312176 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 342192 592650 342812 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 372828 592650 373448 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 403464 592650 404084 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 434100 592650 434720 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 464736 592650 465356 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 495372 592650 495992 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 526008 592650 526628 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 556644 592650 557264 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 587280 592650 587900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 617916 592650 618536 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 648552 592650 649172 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 679188 592650 679808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 198134 17360 198754 139312 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 385262 154448 385882 276400 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 574966 290992 575586 414032 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 198134 154448 198754 276400 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 385262 17360 385882 139312 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 574966 428080 575586 551120 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 198134 291536 198754 413488 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 385262 428624 385882 550576 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 574966 17360 575586 139856 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 198134 428624 198754 550576 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 385262 291536 385882 413488 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 574966 153904 575586 276944 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 198134 565712 198754 687664 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 385262 565712 385882 687664 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 574966 565168 575586 687664 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 4058 148950 582868 149570 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 4058 422990 582868 423610 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 95646330
string GDS_FILE /home/alex/chaos_automaton_Summer_2022/openlane/user_project_wrapper/runs/22_08_12_13_01/results/signoff/user_project_wrapper.magic.gds
string GDS_START 51838014
<< end >>

