VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chaos_subarray
  CLASS BLOCK ;
  FOREIGN chaos_subarray ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN hold
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END hold
  PIN iclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END iclk
  PIN idata
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END idata
  PIN ieast[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 13.640 900.000 14.240 ;
    END
  END ieast[0]
  PIN ieast[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 40.840 900.000 41.440 ;
    END
  END ieast[1]
  PIN ieast[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 68.040 900.000 68.640 ;
    END
  END ieast[2]
  PIN ieast[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 95.240 900.000 95.840 ;
    END
  END ieast[3]
  PIN ieast[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 122.440 900.000 123.040 ;
    END
  END ieast[4]
  PIN ieast[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 149.640 900.000 150.240 ;
    END
  END ieast[5]
  PIN ieast[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 176.840 900.000 177.440 ;
    END
  END ieast[6]
  PIN ieast[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 204.040 900.000 204.640 ;
    END
  END ieast[7]
  PIN ieast[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 231.240 900.000 231.840 ;
    END
  END ieast[8]
  PIN ieast[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 258.440 900.000 259.040 ;
    END
  END ieast[9]
  PIN inorth[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 596.000 873.910 600.000 ;
    END
  END inorth[0]
  PIN inorth[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 596.000 829.290 600.000 ;
    END
  END inorth[1]
  PIN inorth[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 596.000 784.670 600.000 ;
    END
  END inorth[2]
  PIN inorth[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 596.000 740.050 600.000 ;
    END
  END inorth[3]
  PIN inorth[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 596.000 695.430 600.000 ;
    END
  END inorth[4]
  PIN inorth[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 596.000 650.810 600.000 ;
    END
  END inorth[5]
  PIN inorth[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 596.000 606.190 600.000 ;
    END
  END inorth[6]
  PIN inorth[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 596.000 561.570 600.000 ;
    END
  END inorth[7]
  PIN inorth[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 596.000 516.950 600.000 ;
    END
  END inorth[8]
  PIN inorth[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 596.000 472.330 600.000 ;
    END
  END inorth[9]
  PIN isouth[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END isouth[0]
  PIN isouth[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END isouth[1]
  PIN isouth[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END isouth[2]
  PIN isouth[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END isouth[3]
  PIN isouth[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END isouth[4]
  PIN isouth[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END isouth[5]
  PIN isouth[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END isouth[6]
  PIN isouth[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END isouth[7]
  PIN isouth[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END isouth[8]
  PIN isouth[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END isouth[9]
  PIN iwest[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END iwest[0]
  PIN iwest[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END iwest[1]
  PIN iwest[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END iwest[2]
  PIN iwest[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END iwest[3]
  PIN iwest[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END iwest[4]
  PIN iwest[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END iwest[5]
  PIN iwest[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END iwest[6]
  PIN iwest[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END iwest[7]
  PIN iwest[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END iwest[8]
  PIN iwest[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END iwest[9]
  PIN oclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 557.640 900.000 558.240 ;
    END
  END oclk
  PIN odata
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 584.840 900.000 585.440 ;
    END
  END odata
  PIN oeast[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 285.640 900.000 286.240 ;
    END
  END oeast[0]
  PIN oeast[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 312.840 900.000 313.440 ;
    END
  END oeast[1]
  PIN oeast[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 340.040 900.000 340.640 ;
    END
  END oeast[2]
  PIN oeast[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 367.240 900.000 367.840 ;
    END
  END oeast[3]
  PIN oeast[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 394.440 900.000 395.040 ;
    END
  END oeast[4]
  PIN oeast[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 421.640 900.000 422.240 ;
    END
  END oeast[5]
  PIN oeast[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 448.840 900.000 449.440 ;
    END
  END oeast[6]
  PIN oeast[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 476.040 900.000 476.640 ;
    END
  END oeast[7]
  PIN oeast[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 503.240 900.000 503.840 ;
    END
  END oeast[8]
  PIN oeast[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 530.440 900.000 531.040 ;
    END
  END oeast[9]
  PIN onorth[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 596.000 427.710 600.000 ;
    END
  END onorth[0]
  PIN onorth[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 596.000 383.090 600.000 ;
    END
  END onorth[1]
  PIN onorth[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 596.000 338.470 600.000 ;
    END
  END onorth[2]
  PIN onorth[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 596.000 293.850 600.000 ;
    END
  END onorth[3]
  PIN onorth[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 596.000 249.230 600.000 ;
    END
  END onorth[4]
  PIN onorth[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 596.000 204.610 600.000 ;
    END
  END onorth[5]
  PIN onorth[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 596.000 159.990 600.000 ;
    END
  END onorth[6]
  PIN onorth[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 596.000 115.370 600.000 ;
    END
  END onorth[7]
  PIN onorth[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 596.000 70.750 600.000 ;
    END
  END onorth[8]
  PIN onorth[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 596.000 26.130 600.000 ;
    END
  END onorth[9]
  PIN osouth[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END osouth[0]
  PIN osouth[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END osouth[1]
  PIN osouth[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 0.000 591.930 4.000 ;
    END
  END osouth[2]
  PIN osouth[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END osouth[3]
  PIN osouth[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END osouth[4]
  PIN osouth[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 0.000 713.370 4.000 ;
    END
  END osouth[5]
  PIN osouth[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END osouth[6]
  PIN osouth[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 0.000 794.330 4.000 ;
    END
  END osouth[7]
  PIN osouth[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 0.000 834.810 4.000 ;
    END
  END osouth[8]
  PIN osouth[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END osouth[9]
  PIN owest[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END owest[0]
  PIN owest[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END owest[1]
  PIN owest[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END owest[2]
  PIN owest[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END owest[3]
  PIN owest[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END owest[4]
  PIN owest[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END owest[5]
  PIN owest[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END owest[6]
  PIN owest[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END owest[7]
  PIN owest[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END owest[8]
  PIN owest[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END owest[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 894.480 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 894.480 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 894.480 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 894.480 487.870 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 103.320 894.480 104.920 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 256.500 894.480 258.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 409.680 894.480 411.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 562.860 894.480 564.460 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 8.200 894.240 587.760 ;
      LAYER met2 ;
        RECT 6.990 595.720 25.570 596.770 ;
        RECT 26.410 595.720 70.190 596.770 ;
        RECT 71.030 595.720 114.810 596.770 ;
        RECT 115.650 595.720 159.430 596.770 ;
        RECT 160.270 595.720 204.050 596.770 ;
        RECT 204.890 595.720 248.670 596.770 ;
        RECT 249.510 595.720 293.290 596.770 ;
        RECT 294.130 595.720 337.910 596.770 ;
        RECT 338.750 595.720 382.530 596.770 ;
        RECT 383.370 595.720 427.150 596.770 ;
        RECT 427.990 595.720 471.770 596.770 ;
        RECT 472.610 595.720 516.390 596.770 ;
        RECT 517.230 595.720 561.010 596.770 ;
        RECT 561.850 595.720 605.630 596.770 ;
        RECT 606.470 595.720 650.250 596.770 ;
        RECT 651.090 595.720 694.870 596.770 ;
        RECT 695.710 595.720 739.490 596.770 ;
        RECT 740.330 595.720 784.110 596.770 ;
        RECT 784.950 595.720 828.730 596.770 ;
        RECT 829.570 595.720 873.350 596.770 ;
        RECT 874.190 595.720 892.310 596.770 ;
        RECT 6.990 4.280 892.310 595.720 ;
        RECT 6.990 4.000 24.650 4.280 ;
        RECT 25.490 4.000 65.130 4.280 ;
        RECT 65.970 4.000 105.610 4.280 ;
        RECT 106.450 4.000 146.090 4.280 ;
        RECT 146.930 4.000 186.570 4.280 ;
        RECT 187.410 4.000 227.050 4.280 ;
        RECT 227.890 4.000 267.530 4.280 ;
        RECT 268.370 4.000 308.010 4.280 ;
        RECT 308.850 4.000 348.490 4.280 ;
        RECT 349.330 4.000 388.970 4.280 ;
        RECT 389.810 4.000 429.450 4.280 ;
        RECT 430.290 4.000 469.930 4.280 ;
        RECT 470.770 4.000 510.410 4.280 ;
        RECT 511.250 4.000 550.890 4.280 ;
        RECT 551.730 4.000 591.370 4.280 ;
        RECT 592.210 4.000 631.850 4.280 ;
        RECT 632.690 4.000 672.330 4.280 ;
        RECT 673.170 4.000 712.810 4.280 ;
        RECT 713.650 4.000 753.290 4.280 ;
        RECT 754.130 4.000 793.770 4.280 ;
        RECT 794.610 4.000 834.250 4.280 ;
        RECT 835.090 4.000 874.730 4.280 ;
        RECT 875.570 4.000 892.310 4.280 ;
      LAYER met3 ;
        RECT 4.000 585.840 896.000 587.685 ;
        RECT 4.400 584.440 895.600 585.840 ;
        RECT 4.000 558.640 896.000 584.440 ;
        RECT 4.400 557.240 895.600 558.640 ;
        RECT 4.000 531.440 896.000 557.240 ;
        RECT 4.400 530.040 895.600 531.440 ;
        RECT 4.000 504.240 896.000 530.040 ;
        RECT 4.400 502.840 895.600 504.240 ;
        RECT 4.000 477.040 896.000 502.840 ;
        RECT 4.400 475.640 895.600 477.040 ;
        RECT 4.000 449.840 896.000 475.640 ;
        RECT 4.400 448.440 895.600 449.840 ;
        RECT 4.000 422.640 896.000 448.440 ;
        RECT 4.400 421.240 895.600 422.640 ;
        RECT 4.000 395.440 896.000 421.240 ;
        RECT 4.400 394.040 895.600 395.440 ;
        RECT 4.000 368.240 896.000 394.040 ;
        RECT 4.400 366.840 895.600 368.240 ;
        RECT 4.000 341.040 896.000 366.840 ;
        RECT 4.400 339.640 895.600 341.040 ;
        RECT 4.000 313.840 896.000 339.640 ;
        RECT 4.400 312.440 895.600 313.840 ;
        RECT 4.000 286.640 896.000 312.440 ;
        RECT 4.400 285.240 895.600 286.640 ;
        RECT 4.000 259.440 896.000 285.240 ;
        RECT 4.400 258.040 895.600 259.440 ;
        RECT 4.000 232.240 896.000 258.040 ;
        RECT 4.400 230.840 895.600 232.240 ;
        RECT 4.000 205.040 896.000 230.840 ;
        RECT 4.400 203.640 895.600 205.040 ;
        RECT 4.000 177.840 896.000 203.640 ;
        RECT 4.400 176.440 895.600 177.840 ;
        RECT 4.000 150.640 896.000 176.440 ;
        RECT 4.400 149.240 895.600 150.640 ;
        RECT 4.000 123.440 896.000 149.240 ;
        RECT 4.400 122.040 895.600 123.440 ;
        RECT 4.000 96.240 896.000 122.040 ;
        RECT 4.400 94.840 895.600 96.240 ;
        RECT 4.000 69.040 896.000 94.840 ;
        RECT 4.400 67.640 895.600 69.040 ;
        RECT 4.000 41.840 896.000 67.640 ;
        RECT 4.400 40.440 895.600 41.840 ;
        RECT 4.000 14.640 896.000 40.440 ;
        RECT 4.400 13.240 895.600 14.640 ;
        RECT 4.000 10.715 896.000 13.240 ;
      LAYER met4 ;
        RECT 10.415 70.215 20.640 531.585 ;
        RECT 23.040 70.215 97.440 531.585 ;
        RECT 99.840 70.215 174.240 531.585 ;
        RECT 176.640 70.215 251.040 531.585 ;
        RECT 253.440 70.215 327.840 531.585 ;
        RECT 330.240 70.215 404.640 531.585 ;
        RECT 407.040 70.215 481.440 531.585 ;
        RECT 483.840 70.215 558.240 531.585 ;
        RECT 560.640 70.215 635.040 531.585 ;
        RECT 637.440 70.215 711.840 531.585 ;
        RECT 714.240 70.215 788.640 531.585 ;
        RECT 791.040 70.215 865.440 531.585 ;
        RECT 867.840 70.215 889.345 531.585 ;
  END
END chaos_subarray
END LIBRARY

