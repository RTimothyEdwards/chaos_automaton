VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chaos_automaton
  CLASS BLOCK ;
  FOREIGN chaos_automaton ;
  ORIGIN 0.000 0.000 ;
  SIZE 3006.000 BY 3596.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 46.960 3006.000 47.560 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2433.760 3006.000 2434.360 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2672.440 3006.000 2673.040 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2911.120 3006.000 2911.720 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 3149.800 3006.000 3150.400 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 3388.480 3006.000 3389.080 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2950.070 3592.000 2950.350 3596.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2616.110 3592.000 2616.390 3596.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.150 3592.000 2282.430 3596.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.190 3592.000 1948.470 3596.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.230 3592.000 1614.510 3596.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 285.640 3006.000 286.240 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.270 3592.000 1280.550 3596.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 3592.000 946.590 3596.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 3592.000 612.630 3596.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 3592.000 278.670 3596.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3540.120 4.000 3540.720 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3285.120 4.000 3285.720 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3030.120 4.000 3030.720 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2775.120 4.000 2775.720 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2520.120 4.000 2520.720 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2265.120 4.000 2265.720 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 524.320 3006.000 524.920 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2010.120 4.000 2010.720 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1755.120 4.000 1755.720 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1500.120 4.000 1500.720 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1245.120 4.000 1245.720 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.120 4.000 990.720 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.120 4.000 735.720 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 763.000 3006.000 763.600 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1001.680 3006.000 1002.280 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1240.360 3006.000 1240.960 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1479.040 3006.000 1479.640 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1717.720 3006.000 1718.320 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1956.400 3006.000 1957.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2195.080 3006.000 2195.680 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 206.080 3006.000 206.680 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2592.880 3006.000 2593.480 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2831.560 3006.000 2832.160 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 3070.240 3006.000 3070.840 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 3308.920 3006.000 3309.520 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 3547.600 3006.000 3548.200 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.430 3592.000 2727.710 3596.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2393.470 3592.000 2393.750 3596.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.510 3592.000 2059.790 3596.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.550 3592.000 1725.830 3596.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.590 3592.000 1391.870 3596.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 444.760 3006.000 445.360 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.630 3592.000 1057.910 3596.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 3592.000 723.950 3596.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 3592.000 389.990 3596.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 3592.000 56.030 3596.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3370.120 4.000 3370.720 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3115.120 4.000 3115.720 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2860.120 4.000 2860.720 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2605.120 4.000 2605.720 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2350.120 4.000 2350.720 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2095.120 4.000 2095.720 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 683.440 3006.000 684.040 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1840.120 4.000 1840.720 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1585.120 4.000 1585.720 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1330.120 4.000 1330.720 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1075.120 4.000 1075.720 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.120 4.000 820.720 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.120 4.000 565.720 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 922.120 3006.000 922.720 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1160.800 3006.000 1161.400 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1399.480 3006.000 1400.080 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1638.160 3006.000 1638.760 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1876.840 3006.000 1877.440 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2115.520 3006.000 2116.120 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2354.200 3006.000 2354.800 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 126.520 3006.000 127.120 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2513.320 3006.000 2513.920 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2752.000 3006.000 2752.600 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2990.680 3006.000 2991.280 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 3229.360 3006.000 3229.960 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 3468.040 3006.000 3468.640 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2838.750 3592.000 2839.030 3596.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2504.790 3592.000 2505.070 3596.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2170.830 3592.000 2171.110 3596.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1836.870 3592.000 1837.150 3596.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1502.910 3592.000 1503.190 3596.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 365.200 3006.000 365.800 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 3592.000 1169.230 3596.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 3592.000 835.270 3596.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 3592.000 501.310 3596.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 3592.000 167.350 3596.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3455.120 4.000 3455.720 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3200.120 4.000 3200.720 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2945.120 4.000 2945.720 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2690.120 4.000 2690.720 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2435.120 4.000 2435.720 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2180.120 4.000 2180.720 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 603.880 3006.000 604.480 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1925.120 4.000 1925.720 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1670.120 4.000 1670.720 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1415.120 4.000 1415.720 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1160.120 4.000 1160.720 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.120 4.000 905.720 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 842.560 3006.000 843.160 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1081.240 3006.000 1081.840 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1319.920 3006.000 1320.520 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1558.600 3006.000 1559.200 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 1797.280 3006.000 1797.880 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2035.960 3006.000 2036.560 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3002.000 2274.640 3006.000 2275.240 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2962.030 0.000 2962.310 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2968.010 0.000 2968.290 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2973.990 0.000 2974.270 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2459.710 0.000 2459.990 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2477.650 0.000 2477.930 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2495.590 0.000 2495.870 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2513.530 0.000 2513.810 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2531.470 0.000 2531.750 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2549.410 0.000 2549.690 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.350 0.000 2567.630 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.290 0.000 2585.570 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.230 0.000 2603.510 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.170 0.000 2621.450 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 0.000 845.390 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2639.110 0.000 2639.390 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2657.050 0.000 2657.330 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.990 0.000 2675.270 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2692.930 0.000 2693.210 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2710.870 0.000 2711.150 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2728.810 0.000 2729.090 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2746.750 0.000 2747.030 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2764.690 0.000 2764.970 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2782.630 0.000 2782.910 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2800.570 0.000 2800.850 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2818.510 0.000 2818.790 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2836.450 0.000 2836.730 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2854.390 0.000 2854.670 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2872.330 0.000 2872.610 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2890.270 0.000 2890.550 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2908.210 0.000 2908.490 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2926.150 0.000 2926.430 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2944.090 0.000 2944.370 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 0.000 881.270 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.930 0.000 899.210 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.870 0.000 917.150 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 0.000 935.090 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 0.000 953.030 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.690 0.000 970.970 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.570 0.000 1006.850 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.510 0.000 1024.790 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.450 0.000 1042.730 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.390 0.000 1060.670 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.330 0.000 1078.610 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.270 0.000 1096.550 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.150 0.000 1132.430 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 0.000 1150.370 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.030 0.000 1168.310 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.970 0.000 1186.250 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 0.000 701.870 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.910 0.000 1204.190 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.850 0.000 1222.130 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 0.000 1240.070 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.730 0.000 1258.010 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.670 0.000 1275.950 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.610 0.000 1293.890 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.550 0.000 1311.830 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.490 0.000 1329.770 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1347.430 0.000 1347.710 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.370 0.000 1365.650 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 0.000 719.810 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1383.310 0.000 1383.590 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.250 0.000 1401.530 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.190 0.000 1419.470 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.130 0.000 1437.410 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.070 0.000 1455.350 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.010 0.000 1473.290 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 0.000 1491.230 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.890 0.000 1509.170 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.830 0.000 1527.110 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.770 0.000 1545.050 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.710 0.000 1562.990 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.650 0.000 1580.930 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.590 0.000 1598.870 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 0.000 1616.810 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.470 0.000 1634.750 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.410 0.000 1652.690 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.350 0.000 1670.630 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.290 0.000 1688.570 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.230 0.000 1706.510 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.170 0.000 1724.450 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 0.000 755.690 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.110 0.000 1742.390 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.050 0.000 1760.330 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.990 0.000 1778.270 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.930 0.000 1796.210 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1813.870 0.000 1814.150 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1831.810 0.000 1832.090 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.750 0.000 1850.030 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1867.690 0.000 1867.970 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1885.630 0.000 1885.910 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.570 0.000 1903.850 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 0.000 773.630 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1921.510 0.000 1921.790 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1939.450 0.000 1939.730 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.390 0.000 1957.670 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.330 0.000 1975.610 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1993.270 0.000 1993.550 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2011.210 0.000 2011.490 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.150 0.000 2029.430 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.090 0.000 2047.370 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.030 0.000 2065.310 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.970 0.000 2083.250 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 0.000 791.570 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.910 0.000 2101.190 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.850 0.000 2119.130 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.790 0.000 2137.070 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.730 0.000 2155.010 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.670 0.000 2172.950 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.610 0.000 2190.890 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2208.550 0.000 2208.830 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2226.490 0.000 2226.770 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2244.430 0.000 2244.710 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.370 0.000 2262.650 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 0.000 809.510 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2280.310 0.000 2280.590 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2298.250 0.000 2298.530 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2316.190 0.000 2316.470 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.130 0.000 2334.410 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2352.070 0.000 2352.350 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2370.010 0.000 2370.290 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2387.950 0.000 2388.230 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.890 0.000 2406.170 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2423.830 0.000 2424.110 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2441.770 0.000 2442.050 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.170 0.000 827.450 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2465.690 0.000 2465.970 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2483.630 0.000 2483.910 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2501.570 0.000 2501.850 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2519.510 0.000 2519.790 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2537.450 0.000 2537.730 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2555.390 0.000 2555.670 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.330 0.000 2573.610 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.270 0.000 2591.550 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.210 0.000 2609.490 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.150 0.000 2627.430 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2645.090 0.000 2645.370 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2663.030 0.000 2663.310 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.970 0.000 2681.250 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2698.910 0.000 2699.190 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2716.850 0.000 2717.130 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2734.790 0.000 2735.070 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2752.730 0.000 2753.010 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2770.670 0.000 2770.950 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2788.610 0.000 2788.890 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2806.550 0.000 2806.830 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.030 0.000 869.310 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2824.490 0.000 2824.770 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2842.430 0.000 2842.710 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2860.370 0.000 2860.650 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2878.310 0.000 2878.590 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2896.250 0.000 2896.530 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2914.190 0.000 2914.470 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2932.130 0.000 2932.410 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2950.070 0.000 2950.350 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.970 0.000 887.250 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.850 0.000 923.130 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.790 0.000 941.070 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730 0.000 959.010 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 0.000 976.950 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.610 0.000 994.890 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.550 0.000 1012.830 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.430 0.000 1048.710 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 0.000 1066.650 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 0.000 1084.590 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 0.000 1102.530 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.190 0.000 1120.470 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 0.000 1138.410 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.010 0.000 1174.290 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 0.000 1192.230 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.890 0.000 1210.170 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.830 0.000 1228.110 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.770 0.000 1246.050 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.710 0.000 1263.990 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.650 0.000 1281.930 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.590 0.000 1299.870 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.530 0.000 1317.810 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.470 0.000 1335.750 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1353.410 0.000 1353.690 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.350 0.000 1371.630 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 0.000 725.790 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1389.290 0.000 1389.570 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 0.000 1407.510 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.170 0.000 1425.450 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.110 0.000 1443.390 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.050 0.000 1461.330 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.990 0.000 1479.270 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.930 0.000 1497.210 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.870 0.000 1515.150 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 0.000 1533.090 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.750 0.000 1551.030 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 0.000 743.730 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.690 0.000 1568.970 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.630 0.000 1586.910 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.570 0.000 1604.850 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.510 0.000 1622.790 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1640.450 0.000 1640.730 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.390 0.000 1658.670 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1676.330 0.000 1676.610 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.270 0.000 1694.550 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.210 0.000 1712.490 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1730.150 0.000 1730.430 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 0.000 761.670 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.090 0.000 1748.370 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.030 0.000 1766.310 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.970 0.000 1784.250 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.910 0.000 1802.190 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.850 0.000 1820.130 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.790 0.000 1838.070 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1855.730 0.000 1856.010 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1873.670 0.000 1873.950 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1891.610 0.000 1891.890 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.550 0.000 1909.830 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.490 0.000 1927.770 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.430 0.000 1945.710 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1963.370 0.000 1963.650 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.310 0.000 1981.590 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1999.250 0.000 1999.530 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.190 0.000 2017.470 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.130 0.000 2035.410 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.070 0.000 2053.350 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.010 0.000 2071.290 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2088.950 0.000 2089.230 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 0.000 797.550 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.890 0.000 2107.170 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.830 0.000 2125.110 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.770 0.000 2143.050 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.710 0.000 2160.990 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2178.650 0.000 2178.930 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.590 0.000 2196.870 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2214.530 0.000 2214.810 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.470 0.000 2232.750 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2250.410 0.000 2250.690 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.350 0.000 2268.630 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.290 0.000 2286.570 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2304.230 0.000 2304.510 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2322.170 0.000 2322.450 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2340.110 0.000 2340.390 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2358.050 0.000 2358.330 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2375.990 0.000 2376.270 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2393.930 0.000 2394.210 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.870 0.000 2412.150 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2429.810 0.000 2430.090 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2447.750 0.000 2448.030 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 0.000 833.430 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 0.000 677.950 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2471.670 0.000 2471.950 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.610 0.000 2489.890 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2507.550 0.000 2507.830 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2525.490 0.000 2525.770 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2543.430 0.000 2543.710 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2561.370 0.000 2561.650 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.310 0.000 2579.590 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.250 0.000 2597.530 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.190 0.000 2615.470 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2633.130 0.000 2633.410 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.070 0.000 857.350 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2651.070 0.000 2651.350 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2669.010 0.000 2669.290 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2686.950 0.000 2687.230 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2704.890 0.000 2705.170 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2722.830 0.000 2723.110 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2740.770 0.000 2741.050 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2758.710 0.000 2758.990 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2776.650 0.000 2776.930 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2794.590 0.000 2794.870 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2812.530 0.000 2812.810 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2830.470 0.000 2830.750 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2848.410 0.000 2848.690 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2866.350 0.000 2866.630 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2884.290 0.000 2884.570 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2902.230 0.000 2902.510 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2920.170 0.000 2920.450 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2938.110 0.000 2938.390 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2956.050 0.000 2956.330 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.950 0.000 893.230 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 0.000 911.170 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 0.000 929.110 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 0.000 964.990 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 0.000 982.930 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 0.000 1000.870 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.530 0.000 1018.810 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.470 0.000 1036.750 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.410 0.000 1054.690 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.290 0.000 1090.570 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.230 0.000 1108.510 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.170 0.000 1126.450 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.110 0.000 1144.390 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.050 0.000 1162.330 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.990 0.000 1180.270 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 0.000 1198.210 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.870 0.000 1216.150 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.810 0.000 1234.090 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.750 0.000 1252.030 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.690 0.000 1269.970 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.630 0.000 1287.910 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.570 0.000 1305.850 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.450 0.000 1341.730 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.390 0.000 1359.670 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.330 0.000 1377.610 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.270 0.000 1395.550 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.210 0.000 1413.490 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.150 0.000 1431.430 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.030 0.000 1467.310 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.970 0.000 1485.250 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1502.910 0.000 1503.190 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1520.850 0.000 1521.130 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1538.790 0.000 1539.070 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.730 0.000 1557.010 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.670 0.000 1574.950 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.610 0.000 1592.890 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.550 0.000 1610.830 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.490 0.000 1628.770 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.430 0.000 1646.710 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.370 0.000 1664.650 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.310 0.000 1682.590 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 0.000 1700.530 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.190 0.000 1718.470 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.130 0.000 1736.410 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.070 0.000 1754.350 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.010 0.000 1772.290 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1789.950 0.000 1790.230 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1807.890 0.000 1808.170 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.830 0.000 1826.110 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1843.770 0.000 1844.050 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.710 0.000 1861.990 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1879.650 0.000 1879.930 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1897.590 0.000 1897.870 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.530 0.000 1915.810 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.470 0.000 1933.750 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.410 0.000 1951.690 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.350 0.000 1969.630 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.290 0.000 1987.570 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2005.230 0.000 2005.510 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.170 0.000 2023.450 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.110 0.000 2041.390 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.050 0.000 2059.330 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.990 0.000 2077.270 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.930 0.000 2095.210 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.250 0.000 803.530 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.870 0.000 2113.150 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.810 0.000 2131.090 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.750 0.000 2149.030 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.690 0.000 2166.970 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2184.630 0.000 2184.910 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.570 0.000 2202.850 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2220.510 0.000 2220.790 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2238.450 0.000 2238.730 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2256.390 0.000 2256.670 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2274.330 0.000 2274.610 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.270 0.000 2292.550 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2310.210 0.000 2310.490 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.150 0.000 2328.430 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2346.090 0.000 2346.370 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2364.030 0.000 2364.310 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2381.970 0.000 2382.250 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2399.910 0.000 2400.190 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.850 0.000 2418.130 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2435.790 0.000 2436.070 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2453.730 0.000 2454.010 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 0.000 839.410 4.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 3592.560 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 3007.720 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3590.960 3007.720 3592.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 3006.120 3.280 3007.720 3592.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.840 -0.020 30.840 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 166.440 -0.020 184.440 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 166.440 730.000 184.440 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 166.440 1429.000 184.440 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 166.440 2128.000 184.440 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 166.440 2827.000 184.440 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 166.440 3526.000 184.440 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 320.040 -0.020 338.040 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 320.040 730.000 338.040 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 320.040 1429.000 338.040 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 320.040 2128.000 338.040 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 320.040 2827.000 338.040 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 320.040 3526.000 338.040 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.640 -0.020 491.640 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.640 730.000 491.640 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.640 1429.000 491.640 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.640 2128.000 491.640 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.640 2827.000 491.640 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.640 3526.000 491.640 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.240 -0.020 645.240 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.240 730.000 645.240 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.240 1429.000 645.240 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.240 2128.000 645.240 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.240 2827.000 645.240 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.240 3526.000 645.240 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 780.840 -0.020 798.840 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 780.840 730.000 798.840 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 780.840 1429.000 798.840 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 780.840 2128.000 798.840 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 780.840 2827.000 798.840 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 780.840 3526.000 798.840 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 934.440 -0.020 952.440 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 934.440 730.000 952.440 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 934.440 1429.000 952.440 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 934.440 2128.000 952.440 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 934.440 2827.000 952.440 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 934.440 3526.000 952.440 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.040 -0.020 1106.040 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.040 730.000 1106.040 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.040 1429.000 1106.040 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.040 2128.000 1106.040 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.040 2827.000 1106.040 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.040 3526.000 1106.040 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1241.640 -0.020 1259.640 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1241.640 730.000 1259.640 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1241.640 1429.000 1259.640 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1241.640 2128.000 1259.640 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1241.640 2827.000 1259.640 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1241.640 3526.000 1259.640 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.240 -0.020 1413.240 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.240 730.000 1413.240 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.240 1429.000 1413.240 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.240 2128.000 1413.240 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.240 2827.000 1413.240 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.240 3526.000 1413.240 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.840 -0.020 1566.840 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.840 730.000 1566.840 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.840 1429.000 1566.840 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.840 2128.000 1566.840 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.840 2827.000 1566.840 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.840 3526.000 1566.840 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1702.440 -0.020 1720.440 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1702.440 730.000 1720.440 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1702.440 1429.000 1720.440 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1702.440 2128.000 1720.440 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1702.440 2827.000 1720.440 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1702.440 3526.000 1720.440 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1856.040 -0.020 1874.040 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1856.040 730.000 1874.040 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1856.040 1429.000 1874.040 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1856.040 2128.000 1874.040 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1856.040 2827.000 1874.040 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1856.040 3526.000 1874.040 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2009.640 -0.020 2027.640 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2009.640 730.000 2027.640 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2009.640 1429.000 2027.640 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2009.640 2128.000 2027.640 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2009.640 2827.000 2027.640 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2009.640 3526.000 2027.640 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2163.240 -0.020 2181.240 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2163.240 730.000 2181.240 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2163.240 1429.000 2181.240 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2163.240 2128.000 2181.240 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2163.240 2827.000 2181.240 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2163.240 3526.000 2181.240 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2316.840 -0.020 2334.840 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2316.840 730.000 2334.840 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2316.840 1429.000 2334.840 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2316.840 2128.000 2334.840 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2316.840 2827.000 2334.840 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2316.840 3526.000 2334.840 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2470.440 -0.020 2488.440 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2470.440 730.000 2488.440 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2470.440 1429.000 2488.440 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2470.440 2128.000 2488.440 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2470.440 2827.000 2488.440 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2470.440 3526.000 2488.440 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2624.040 -0.020 2642.040 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2624.040 730.000 2642.040 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2624.040 1429.000 2642.040 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2624.040 2128.000 2642.040 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2624.040 2827.000 2642.040 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2624.040 3526.000 2642.040 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2777.640 -0.020 2795.640 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2777.640 730.000 2795.640 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2777.640 1429.000 2795.640 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2777.640 2128.000 2795.640 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2777.640 2827.000 2795.640 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2777.640 3526.000 2795.640 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.240 -0.020 2949.240 3595.860 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 19.030 3011.020 36.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 172.210 3011.020 189.210 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 325.390 3011.020 342.390 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 478.570 3011.020 495.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 631.750 3011.020 648.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 784.930 3011.020 801.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 938.110 3011.020 955.110 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1091.290 3011.020 1108.290 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1244.470 3011.020 1261.470 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1397.650 3011.020 1414.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1550.830 3011.020 1567.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1704.010 3011.020 1721.010 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1857.190 3011.020 1874.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2010.370 3011.020 2027.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2163.550 3011.020 2180.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2316.730 3011.020 2333.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2469.910 3011.020 2486.910 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2623.090 3011.020 2640.090 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2776.270 3011.020 2793.270 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2929.450 3011.020 2946.450 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 3082.630 3011.020 3099.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 3235.810 3011.020 3252.810 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 3388.990 3011.020 3405.990 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 3542.170 3011.020 3559.170 ;
    END
    PORT
      LAYER met4 ;
        RECT 1030.040 807.600 1039.040 1433.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1970.280 1503.920 1979.280 2132.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1030.040 105.840 1039.040 731.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1970.280 2202.960 1979.280 2845.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1030.040 2205.680 1039.040 2845.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1970.280 105.840 1979.280 734.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1030.040 1503.920 1039.040 2130.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1970.280 804.880 1979.280 1433.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1030.040 2902.000 1039.040 3528.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1970.280 2902.000 1979.280 3530.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 12.840 1441.600 2949.240 1458.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 12.840 2828.800 2949.240 2845.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 3595.860 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 3011.020 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 3594.260 3011.020 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 3009.420 -0.020 3011.020 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.640 -0.020 107.640 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.640 730.000 107.640 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.640 1429.000 107.640 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.640 2128.000 107.640 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.640 2827.000 107.640 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.640 3526.000 107.640 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.240 -0.020 261.240 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.240 730.000 261.240 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.240 1429.000 261.240 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.240 2128.000 261.240 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.240 2827.000 261.240 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.240 3526.000 261.240 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.840 -0.020 414.840 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.840 730.000 414.840 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.840 1429.000 414.840 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.840 2128.000 414.840 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.840 2827.000 414.840 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.840 3526.000 414.840 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 550.440 -0.020 568.440 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 550.440 730.000 568.440 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 550.440 1429.000 568.440 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 550.440 2128.000 568.440 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 550.440 2827.000 568.440 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 550.440 3526.000 568.440 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.040 -0.020 722.040 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.040 730.000 722.040 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.040 1429.000 722.040 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.040 2128.000 722.040 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.040 2827.000 722.040 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.040 3526.000 722.040 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 857.640 -0.020 875.640 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 857.640 730.000 875.640 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 857.640 1429.000 875.640 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 857.640 2128.000 875.640 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 857.640 2827.000 875.640 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 857.640 3526.000 875.640 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.240 -0.020 1029.240 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.840 -0.020 1182.840 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.840 730.000 1182.840 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.840 1429.000 1182.840 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.840 2128.000 1182.840 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.840 2827.000 1182.840 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.840 3526.000 1182.840 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1318.440 -0.020 1336.440 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1318.440 730.000 1336.440 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1318.440 1429.000 1336.440 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1318.440 2128.000 1336.440 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1318.440 2827.000 1336.440 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1318.440 3526.000 1336.440 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1472.040 -0.020 1490.040 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1472.040 730.000 1490.040 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1472.040 1429.000 1490.040 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1472.040 2128.000 1490.040 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1472.040 2827.000 1490.040 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1472.040 3526.000 1490.040 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1625.640 -0.020 1643.640 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1625.640 730.000 1643.640 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1625.640 1429.000 1643.640 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1625.640 2128.000 1643.640 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1625.640 2827.000 1643.640 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1625.640 3526.000 1643.640 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1779.240 -0.020 1797.240 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1779.240 730.000 1797.240 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1779.240 1429.000 1797.240 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1779.240 2128.000 1797.240 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1779.240 2827.000 1797.240 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1779.240 3526.000 1797.240 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1932.840 -0.020 1950.840 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1932.840 730.000 1950.840 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1932.840 1429.000 1950.840 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1932.840 2128.000 1950.840 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1932.840 2827.000 1950.840 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1932.840 3526.000 1950.840 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.440 -0.020 2104.440 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.440 730.000 2104.440 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.440 1429.000 2104.440 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.440 2128.000 2104.440 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.440 2827.000 2104.440 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.440 3526.000 2104.440 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2240.040 -0.020 2258.040 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2240.040 730.000 2258.040 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2240.040 1429.000 2258.040 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2240.040 2128.000 2258.040 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2240.040 2827.000 2258.040 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2240.040 3526.000 2258.040 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2393.640 -0.020 2411.640 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2393.640 730.000 2411.640 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2393.640 1429.000 2411.640 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2393.640 2128.000 2411.640 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2393.640 2827.000 2411.640 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2393.640 3526.000 2411.640 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.240 -0.020 2565.240 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.240 730.000 2565.240 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.240 1429.000 2565.240 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.240 2128.000 2565.240 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.240 2827.000 2565.240 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.240 3526.000 2565.240 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.840 -0.020 2718.840 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.840 730.000 2718.840 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.840 1429.000 2718.840 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.840 2128.000 2718.840 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.840 2827.000 2718.840 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.840 3526.000 2718.840 3595.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.440 -0.020 2872.440 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.440 730.000 2872.440 809.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.440 1429.000 2872.440 1508.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.440 2128.000 2872.440 2207.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.440 2827.000 2872.440 2906.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.440 3526.000 2872.440 3595.860 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 95.620 3011.020 112.620 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 248.800 3011.020 265.800 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 401.980 3011.020 418.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 555.160 3011.020 572.160 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 708.340 3011.020 725.340 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 861.520 3011.020 878.520 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1014.700 3011.020 1031.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1167.880 3011.020 1184.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1321.060 3011.020 1338.060 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1474.240 3011.020 1491.240 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1627.420 3011.020 1644.420 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1780.600 3011.020 1797.600 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1933.780 3011.020 1950.780 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2086.960 3011.020 2103.960 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2240.140 3011.020 2257.140 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2393.320 3011.020 2410.320 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2546.500 3011.020 2563.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2699.680 3011.020 2716.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 2852.860 3011.020 2869.860 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 3006.040 3011.020 3023.040 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 3159.220 3011.020 3176.220 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 3312.400 3011.020 3329.400 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 3465.580 3011.020 3482.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.380 95.620 56.380 734.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1980.400 1503.920 1989.400 2132.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2970.420 2202.960 2988.420 2829.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.380 804.880 56.380 1430.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1980.400 2202.960 1989.400 2831.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2970.420 1506.640 2988.420 2132.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.380 1506.640 56.380 2132.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1980.400 95.620 1989.400 734.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 2970.420 804.880 2988.420 1430.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.380 2202.960 56.380 2829.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1980.400 804.880 1989.400 1433.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2970.420 95.620 2988.420 734.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.380 2904.720 56.380 3530.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1980.400 2902.000 1989.400 3530.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2970.420 2904.720 2988.420 3530.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 761.600 3000.360 778.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2138.600 3000.360 2155.600 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 0.000 558.350 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 0.000 576.290 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 0.000 630.110 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 0.000 648.050 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 0.000 510.510 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 0.000 600.210 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 0.000 480.610 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 0.000 498.550 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 0.000 642.070 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 0.000 660.010 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 3000.120 3585.045 ;
      LAYER met1 ;
        RECT 5.520 1.400 3000.120 3586.620 ;
      LAYER met2 ;
        RECT 6.990 3591.720 55.470 3592.000 ;
        RECT 56.310 3591.720 166.790 3592.000 ;
        RECT 167.630 3591.720 278.110 3592.000 ;
        RECT 278.950 3591.720 389.430 3592.000 ;
        RECT 390.270 3591.720 500.750 3592.000 ;
        RECT 501.590 3591.720 612.070 3592.000 ;
        RECT 612.910 3591.720 723.390 3592.000 ;
        RECT 724.230 3591.720 834.710 3592.000 ;
        RECT 835.550 3591.720 946.030 3592.000 ;
        RECT 946.870 3591.720 1057.350 3592.000 ;
        RECT 1058.190 3591.720 1168.670 3592.000 ;
        RECT 1169.510 3591.720 1279.990 3592.000 ;
        RECT 1280.830 3591.720 1391.310 3592.000 ;
        RECT 1392.150 3591.720 1502.630 3592.000 ;
        RECT 1503.470 3591.720 1613.950 3592.000 ;
        RECT 1614.790 3591.720 1725.270 3592.000 ;
        RECT 1726.110 3591.720 1836.590 3592.000 ;
        RECT 1837.430 3591.720 1947.910 3592.000 ;
        RECT 1948.750 3591.720 2059.230 3592.000 ;
        RECT 2060.070 3591.720 2170.550 3592.000 ;
        RECT 2171.390 3591.720 2281.870 3592.000 ;
        RECT 2282.710 3591.720 2393.190 3592.000 ;
        RECT 2394.030 3591.720 2504.510 3592.000 ;
        RECT 2505.350 3591.720 2615.830 3592.000 ;
        RECT 2616.670 3591.720 2727.150 3592.000 ;
        RECT 2727.990 3591.720 2838.470 3592.000 ;
        RECT 2839.310 3591.720 2949.790 3592.000 ;
        RECT 2950.630 3591.720 2997.730 3592.000 ;
        RECT 6.990 4.280 2997.730 3591.720 ;
        RECT 6.990 0.835 31.550 4.280 ;
        RECT 32.390 0.835 37.530 4.280 ;
        RECT 38.370 0.835 43.510 4.280 ;
        RECT 44.350 0.835 49.490 4.280 ;
        RECT 50.330 0.835 55.470 4.280 ;
        RECT 56.310 0.835 61.450 4.280 ;
        RECT 62.290 0.835 67.430 4.280 ;
        RECT 68.270 0.835 73.410 4.280 ;
        RECT 74.250 0.835 79.390 4.280 ;
        RECT 80.230 0.835 85.370 4.280 ;
        RECT 86.210 0.835 91.350 4.280 ;
        RECT 92.190 0.835 97.330 4.280 ;
        RECT 98.170 0.835 103.310 4.280 ;
        RECT 104.150 0.835 109.290 4.280 ;
        RECT 110.130 0.835 115.270 4.280 ;
        RECT 116.110 0.835 121.250 4.280 ;
        RECT 122.090 0.835 127.230 4.280 ;
        RECT 128.070 0.835 133.210 4.280 ;
        RECT 134.050 0.835 139.190 4.280 ;
        RECT 140.030 0.835 145.170 4.280 ;
        RECT 146.010 0.835 151.150 4.280 ;
        RECT 151.990 0.835 157.130 4.280 ;
        RECT 157.970 0.835 163.110 4.280 ;
        RECT 163.950 0.835 169.090 4.280 ;
        RECT 169.930 0.835 175.070 4.280 ;
        RECT 175.910 0.835 181.050 4.280 ;
        RECT 181.890 0.835 187.030 4.280 ;
        RECT 187.870 0.835 193.010 4.280 ;
        RECT 193.850 0.835 198.990 4.280 ;
        RECT 199.830 0.835 204.970 4.280 ;
        RECT 205.810 0.835 210.950 4.280 ;
        RECT 211.790 0.835 216.930 4.280 ;
        RECT 217.770 0.835 222.910 4.280 ;
        RECT 223.750 0.835 228.890 4.280 ;
        RECT 229.730 0.835 234.870 4.280 ;
        RECT 235.710 0.835 240.850 4.280 ;
        RECT 241.690 0.835 246.830 4.280 ;
        RECT 247.670 0.835 252.810 4.280 ;
        RECT 253.650 0.835 258.790 4.280 ;
        RECT 259.630 0.835 264.770 4.280 ;
        RECT 265.610 0.835 270.750 4.280 ;
        RECT 271.590 0.835 276.730 4.280 ;
        RECT 277.570 0.835 282.710 4.280 ;
        RECT 283.550 0.835 288.690 4.280 ;
        RECT 289.530 0.835 294.670 4.280 ;
        RECT 295.510 0.835 300.650 4.280 ;
        RECT 301.490 0.835 306.630 4.280 ;
        RECT 307.470 0.835 312.610 4.280 ;
        RECT 313.450 0.835 318.590 4.280 ;
        RECT 319.430 0.835 324.570 4.280 ;
        RECT 325.410 0.835 330.550 4.280 ;
        RECT 331.390 0.835 336.530 4.280 ;
        RECT 337.370 0.835 342.510 4.280 ;
        RECT 343.350 0.835 348.490 4.280 ;
        RECT 349.330 0.835 354.470 4.280 ;
        RECT 355.310 0.835 360.450 4.280 ;
        RECT 361.290 0.835 366.430 4.280 ;
        RECT 367.270 0.835 372.410 4.280 ;
        RECT 373.250 0.835 378.390 4.280 ;
        RECT 379.230 0.835 384.370 4.280 ;
        RECT 385.210 0.835 390.350 4.280 ;
        RECT 391.190 0.835 396.330 4.280 ;
        RECT 397.170 0.835 402.310 4.280 ;
        RECT 403.150 0.835 408.290 4.280 ;
        RECT 409.130 0.835 414.270 4.280 ;
        RECT 415.110 0.835 420.250 4.280 ;
        RECT 421.090 0.835 426.230 4.280 ;
        RECT 427.070 0.835 432.210 4.280 ;
        RECT 433.050 0.835 438.190 4.280 ;
        RECT 439.030 0.835 444.170 4.280 ;
        RECT 445.010 0.835 450.150 4.280 ;
        RECT 450.990 0.835 456.130 4.280 ;
        RECT 456.970 0.835 462.110 4.280 ;
        RECT 462.950 0.835 468.090 4.280 ;
        RECT 468.930 0.835 474.070 4.280 ;
        RECT 474.910 0.835 480.050 4.280 ;
        RECT 480.890 0.835 486.030 4.280 ;
        RECT 486.870 0.835 492.010 4.280 ;
        RECT 492.850 0.835 497.990 4.280 ;
        RECT 498.830 0.835 503.970 4.280 ;
        RECT 504.810 0.835 509.950 4.280 ;
        RECT 510.790 0.835 515.930 4.280 ;
        RECT 516.770 0.835 521.910 4.280 ;
        RECT 522.750 0.835 527.890 4.280 ;
        RECT 528.730 0.835 533.870 4.280 ;
        RECT 534.710 0.835 539.850 4.280 ;
        RECT 540.690 0.835 545.830 4.280 ;
        RECT 546.670 0.835 551.810 4.280 ;
        RECT 552.650 0.835 557.790 4.280 ;
        RECT 558.630 0.835 563.770 4.280 ;
        RECT 564.610 0.835 569.750 4.280 ;
        RECT 570.590 0.835 575.730 4.280 ;
        RECT 576.570 0.835 581.710 4.280 ;
        RECT 582.550 0.835 587.690 4.280 ;
        RECT 588.530 0.835 593.670 4.280 ;
        RECT 594.510 0.835 599.650 4.280 ;
        RECT 600.490 0.835 605.630 4.280 ;
        RECT 606.470 0.835 611.610 4.280 ;
        RECT 612.450 0.835 617.590 4.280 ;
        RECT 618.430 0.835 623.570 4.280 ;
        RECT 624.410 0.835 629.550 4.280 ;
        RECT 630.390 0.835 635.530 4.280 ;
        RECT 636.370 0.835 641.510 4.280 ;
        RECT 642.350 0.835 647.490 4.280 ;
        RECT 648.330 0.835 653.470 4.280 ;
        RECT 654.310 0.835 659.450 4.280 ;
        RECT 660.290 0.835 665.430 4.280 ;
        RECT 666.270 0.835 671.410 4.280 ;
        RECT 672.250 0.835 677.390 4.280 ;
        RECT 678.230 0.835 683.370 4.280 ;
        RECT 684.210 0.835 689.350 4.280 ;
        RECT 690.190 0.835 695.330 4.280 ;
        RECT 696.170 0.835 701.310 4.280 ;
        RECT 702.150 0.835 707.290 4.280 ;
        RECT 708.130 0.835 713.270 4.280 ;
        RECT 714.110 0.835 719.250 4.280 ;
        RECT 720.090 0.835 725.230 4.280 ;
        RECT 726.070 0.835 731.210 4.280 ;
        RECT 732.050 0.835 737.190 4.280 ;
        RECT 738.030 0.835 743.170 4.280 ;
        RECT 744.010 0.835 749.150 4.280 ;
        RECT 749.990 0.835 755.130 4.280 ;
        RECT 755.970 0.835 761.110 4.280 ;
        RECT 761.950 0.835 767.090 4.280 ;
        RECT 767.930 0.835 773.070 4.280 ;
        RECT 773.910 0.835 779.050 4.280 ;
        RECT 779.890 0.835 785.030 4.280 ;
        RECT 785.870 0.835 791.010 4.280 ;
        RECT 791.850 0.835 796.990 4.280 ;
        RECT 797.830 0.835 802.970 4.280 ;
        RECT 803.810 0.835 808.950 4.280 ;
        RECT 809.790 0.835 814.930 4.280 ;
        RECT 815.770 0.835 820.910 4.280 ;
        RECT 821.750 0.835 826.890 4.280 ;
        RECT 827.730 0.835 832.870 4.280 ;
        RECT 833.710 0.835 838.850 4.280 ;
        RECT 839.690 0.835 844.830 4.280 ;
        RECT 845.670 0.835 850.810 4.280 ;
        RECT 851.650 0.835 856.790 4.280 ;
        RECT 857.630 0.835 862.770 4.280 ;
        RECT 863.610 0.835 868.750 4.280 ;
        RECT 869.590 0.835 874.730 4.280 ;
        RECT 875.570 0.835 880.710 4.280 ;
        RECT 881.550 0.835 886.690 4.280 ;
        RECT 887.530 0.835 892.670 4.280 ;
        RECT 893.510 0.835 898.650 4.280 ;
        RECT 899.490 0.835 904.630 4.280 ;
        RECT 905.470 0.835 910.610 4.280 ;
        RECT 911.450 0.835 916.590 4.280 ;
        RECT 917.430 0.835 922.570 4.280 ;
        RECT 923.410 0.835 928.550 4.280 ;
        RECT 929.390 0.835 934.530 4.280 ;
        RECT 935.370 0.835 940.510 4.280 ;
        RECT 941.350 0.835 946.490 4.280 ;
        RECT 947.330 0.835 952.470 4.280 ;
        RECT 953.310 0.835 958.450 4.280 ;
        RECT 959.290 0.835 964.430 4.280 ;
        RECT 965.270 0.835 970.410 4.280 ;
        RECT 971.250 0.835 976.390 4.280 ;
        RECT 977.230 0.835 982.370 4.280 ;
        RECT 983.210 0.835 988.350 4.280 ;
        RECT 989.190 0.835 994.330 4.280 ;
        RECT 995.170 0.835 1000.310 4.280 ;
        RECT 1001.150 0.835 1006.290 4.280 ;
        RECT 1007.130 0.835 1012.270 4.280 ;
        RECT 1013.110 0.835 1018.250 4.280 ;
        RECT 1019.090 0.835 1024.230 4.280 ;
        RECT 1025.070 0.835 1030.210 4.280 ;
        RECT 1031.050 0.835 1036.190 4.280 ;
        RECT 1037.030 0.835 1042.170 4.280 ;
        RECT 1043.010 0.835 1048.150 4.280 ;
        RECT 1048.990 0.835 1054.130 4.280 ;
        RECT 1054.970 0.835 1060.110 4.280 ;
        RECT 1060.950 0.835 1066.090 4.280 ;
        RECT 1066.930 0.835 1072.070 4.280 ;
        RECT 1072.910 0.835 1078.050 4.280 ;
        RECT 1078.890 0.835 1084.030 4.280 ;
        RECT 1084.870 0.835 1090.010 4.280 ;
        RECT 1090.850 0.835 1095.990 4.280 ;
        RECT 1096.830 0.835 1101.970 4.280 ;
        RECT 1102.810 0.835 1107.950 4.280 ;
        RECT 1108.790 0.835 1113.930 4.280 ;
        RECT 1114.770 0.835 1119.910 4.280 ;
        RECT 1120.750 0.835 1125.890 4.280 ;
        RECT 1126.730 0.835 1131.870 4.280 ;
        RECT 1132.710 0.835 1137.850 4.280 ;
        RECT 1138.690 0.835 1143.830 4.280 ;
        RECT 1144.670 0.835 1149.810 4.280 ;
        RECT 1150.650 0.835 1155.790 4.280 ;
        RECT 1156.630 0.835 1161.770 4.280 ;
        RECT 1162.610 0.835 1167.750 4.280 ;
        RECT 1168.590 0.835 1173.730 4.280 ;
        RECT 1174.570 0.835 1179.710 4.280 ;
        RECT 1180.550 0.835 1185.690 4.280 ;
        RECT 1186.530 0.835 1191.670 4.280 ;
        RECT 1192.510 0.835 1197.650 4.280 ;
        RECT 1198.490 0.835 1203.630 4.280 ;
        RECT 1204.470 0.835 1209.610 4.280 ;
        RECT 1210.450 0.835 1215.590 4.280 ;
        RECT 1216.430 0.835 1221.570 4.280 ;
        RECT 1222.410 0.835 1227.550 4.280 ;
        RECT 1228.390 0.835 1233.530 4.280 ;
        RECT 1234.370 0.835 1239.510 4.280 ;
        RECT 1240.350 0.835 1245.490 4.280 ;
        RECT 1246.330 0.835 1251.470 4.280 ;
        RECT 1252.310 0.835 1257.450 4.280 ;
        RECT 1258.290 0.835 1263.430 4.280 ;
        RECT 1264.270 0.835 1269.410 4.280 ;
        RECT 1270.250 0.835 1275.390 4.280 ;
        RECT 1276.230 0.835 1281.370 4.280 ;
        RECT 1282.210 0.835 1287.350 4.280 ;
        RECT 1288.190 0.835 1293.330 4.280 ;
        RECT 1294.170 0.835 1299.310 4.280 ;
        RECT 1300.150 0.835 1305.290 4.280 ;
        RECT 1306.130 0.835 1311.270 4.280 ;
        RECT 1312.110 0.835 1317.250 4.280 ;
        RECT 1318.090 0.835 1323.230 4.280 ;
        RECT 1324.070 0.835 1329.210 4.280 ;
        RECT 1330.050 0.835 1335.190 4.280 ;
        RECT 1336.030 0.835 1341.170 4.280 ;
        RECT 1342.010 0.835 1347.150 4.280 ;
        RECT 1347.990 0.835 1353.130 4.280 ;
        RECT 1353.970 0.835 1359.110 4.280 ;
        RECT 1359.950 0.835 1365.090 4.280 ;
        RECT 1365.930 0.835 1371.070 4.280 ;
        RECT 1371.910 0.835 1377.050 4.280 ;
        RECT 1377.890 0.835 1383.030 4.280 ;
        RECT 1383.870 0.835 1389.010 4.280 ;
        RECT 1389.850 0.835 1394.990 4.280 ;
        RECT 1395.830 0.835 1400.970 4.280 ;
        RECT 1401.810 0.835 1406.950 4.280 ;
        RECT 1407.790 0.835 1412.930 4.280 ;
        RECT 1413.770 0.835 1418.910 4.280 ;
        RECT 1419.750 0.835 1424.890 4.280 ;
        RECT 1425.730 0.835 1430.870 4.280 ;
        RECT 1431.710 0.835 1436.850 4.280 ;
        RECT 1437.690 0.835 1442.830 4.280 ;
        RECT 1443.670 0.835 1448.810 4.280 ;
        RECT 1449.650 0.835 1454.790 4.280 ;
        RECT 1455.630 0.835 1460.770 4.280 ;
        RECT 1461.610 0.835 1466.750 4.280 ;
        RECT 1467.590 0.835 1472.730 4.280 ;
        RECT 1473.570 0.835 1478.710 4.280 ;
        RECT 1479.550 0.835 1484.690 4.280 ;
        RECT 1485.530 0.835 1490.670 4.280 ;
        RECT 1491.510 0.835 1496.650 4.280 ;
        RECT 1497.490 0.835 1502.630 4.280 ;
        RECT 1503.470 0.835 1508.610 4.280 ;
        RECT 1509.450 0.835 1514.590 4.280 ;
        RECT 1515.430 0.835 1520.570 4.280 ;
        RECT 1521.410 0.835 1526.550 4.280 ;
        RECT 1527.390 0.835 1532.530 4.280 ;
        RECT 1533.370 0.835 1538.510 4.280 ;
        RECT 1539.350 0.835 1544.490 4.280 ;
        RECT 1545.330 0.835 1550.470 4.280 ;
        RECT 1551.310 0.835 1556.450 4.280 ;
        RECT 1557.290 0.835 1562.430 4.280 ;
        RECT 1563.270 0.835 1568.410 4.280 ;
        RECT 1569.250 0.835 1574.390 4.280 ;
        RECT 1575.230 0.835 1580.370 4.280 ;
        RECT 1581.210 0.835 1586.350 4.280 ;
        RECT 1587.190 0.835 1592.330 4.280 ;
        RECT 1593.170 0.835 1598.310 4.280 ;
        RECT 1599.150 0.835 1604.290 4.280 ;
        RECT 1605.130 0.835 1610.270 4.280 ;
        RECT 1611.110 0.835 1616.250 4.280 ;
        RECT 1617.090 0.835 1622.230 4.280 ;
        RECT 1623.070 0.835 1628.210 4.280 ;
        RECT 1629.050 0.835 1634.190 4.280 ;
        RECT 1635.030 0.835 1640.170 4.280 ;
        RECT 1641.010 0.835 1646.150 4.280 ;
        RECT 1646.990 0.835 1652.130 4.280 ;
        RECT 1652.970 0.835 1658.110 4.280 ;
        RECT 1658.950 0.835 1664.090 4.280 ;
        RECT 1664.930 0.835 1670.070 4.280 ;
        RECT 1670.910 0.835 1676.050 4.280 ;
        RECT 1676.890 0.835 1682.030 4.280 ;
        RECT 1682.870 0.835 1688.010 4.280 ;
        RECT 1688.850 0.835 1693.990 4.280 ;
        RECT 1694.830 0.835 1699.970 4.280 ;
        RECT 1700.810 0.835 1705.950 4.280 ;
        RECT 1706.790 0.835 1711.930 4.280 ;
        RECT 1712.770 0.835 1717.910 4.280 ;
        RECT 1718.750 0.835 1723.890 4.280 ;
        RECT 1724.730 0.835 1729.870 4.280 ;
        RECT 1730.710 0.835 1735.850 4.280 ;
        RECT 1736.690 0.835 1741.830 4.280 ;
        RECT 1742.670 0.835 1747.810 4.280 ;
        RECT 1748.650 0.835 1753.790 4.280 ;
        RECT 1754.630 0.835 1759.770 4.280 ;
        RECT 1760.610 0.835 1765.750 4.280 ;
        RECT 1766.590 0.835 1771.730 4.280 ;
        RECT 1772.570 0.835 1777.710 4.280 ;
        RECT 1778.550 0.835 1783.690 4.280 ;
        RECT 1784.530 0.835 1789.670 4.280 ;
        RECT 1790.510 0.835 1795.650 4.280 ;
        RECT 1796.490 0.835 1801.630 4.280 ;
        RECT 1802.470 0.835 1807.610 4.280 ;
        RECT 1808.450 0.835 1813.590 4.280 ;
        RECT 1814.430 0.835 1819.570 4.280 ;
        RECT 1820.410 0.835 1825.550 4.280 ;
        RECT 1826.390 0.835 1831.530 4.280 ;
        RECT 1832.370 0.835 1837.510 4.280 ;
        RECT 1838.350 0.835 1843.490 4.280 ;
        RECT 1844.330 0.835 1849.470 4.280 ;
        RECT 1850.310 0.835 1855.450 4.280 ;
        RECT 1856.290 0.835 1861.430 4.280 ;
        RECT 1862.270 0.835 1867.410 4.280 ;
        RECT 1868.250 0.835 1873.390 4.280 ;
        RECT 1874.230 0.835 1879.370 4.280 ;
        RECT 1880.210 0.835 1885.350 4.280 ;
        RECT 1886.190 0.835 1891.330 4.280 ;
        RECT 1892.170 0.835 1897.310 4.280 ;
        RECT 1898.150 0.835 1903.290 4.280 ;
        RECT 1904.130 0.835 1909.270 4.280 ;
        RECT 1910.110 0.835 1915.250 4.280 ;
        RECT 1916.090 0.835 1921.230 4.280 ;
        RECT 1922.070 0.835 1927.210 4.280 ;
        RECT 1928.050 0.835 1933.190 4.280 ;
        RECT 1934.030 0.835 1939.170 4.280 ;
        RECT 1940.010 0.835 1945.150 4.280 ;
        RECT 1945.990 0.835 1951.130 4.280 ;
        RECT 1951.970 0.835 1957.110 4.280 ;
        RECT 1957.950 0.835 1963.090 4.280 ;
        RECT 1963.930 0.835 1969.070 4.280 ;
        RECT 1969.910 0.835 1975.050 4.280 ;
        RECT 1975.890 0.835 1981.030 4.280 ;
        RECT 1981.870 0.835 1987.010 4.280 ;
        RECT 1987.850 0.835 1992.990 4.280 ;
        RECT 1993.830 0.835 1998.970 4.280 ;
        RECT 1999.810 0.835 2004.950 4.280 ;
        RECT 2005.790 0.835 2010.930 4.280 ;
        RECT 2011.770 0.835 2016.910 4.280 ;
        RECT 2017.750 0.835 2022.890 4.280 ;
        RECT 2023.730 0.835 2028.870 4.280 ;
        RECT 2029.710 0.835 2034.850 4.280 ;
        RECT 2035.690 0.835 2040.830 4.280 ;
        RECT 2041.670 0.835 2046.810 4.280 ;
        RECT 2047.650 0.835 2052.790 4.280 ;
        RECT 2053.630 0.835 2058.770 4.280 ;
        RECT 2059.610 0.835 2064.750 4.280 ;
        RECT 2065.590 0.835 2070.730 4.280 ;
        RECT 2071.570 0.835 2076.710 4.280 ;
        RECT 2077.550 0.835 2082.690 4.280 ;
        RECT 2083.530 0.835 2088.670 4.280 ;
        RECT 2089.510 0.835 2094.650 4.280 ;
        RECT 2095.490 0.835 2100.630 4.280 ;
        RECT 2101.470 0.835 2106.610 4.280 ;
        RECT 2107.450 0.835 2112.590 4.280 ;
        RECT 2113.430 0.835 2118.570 4.280 ;
        RECT 2119.410 0.835 2124.550 4.280 ;
        RECT 2125.390 0.835 2130.530 4.280 ;
        RECT 2131.370 0.835 2136.510 4.280 ;
        RECT 2137.350 0.835 2142.490 4.280 ;
        RECT 2143.330 0.835 2148.470 4.280 ;
        RECT 2149.310 0.835 2154.450 4.280 ;
        RECT 2155.290 0.835 2160.430 4.280 ;
        RECT 2161.270 0.835 2166.410 4.280 ;
        RECT 2167.250 0.835 2172.390 4.280 ;
        RECT 2173.230 0.835 2178.370 4.280 ;
        RECT 2179.210 0.835 2184.350 4.280 ;
        RECT 2185.190 0.835 2190.330 4.280 ;
        RECT 2191.170 0.835 2196.310 4.280 ;
        RECT 2197.150 0.835 2202.290 4.280 ;
        RECT 2203.130 0.835 2208.270 4.280 ;
        RECT 2209.110 0.835 2214.250 4.280 ;
        RECT 2215.090 0.835 2220.230 4.280 ;
        RECT 2221.070 0.835 2226.210 4.280 ;
        RECT 2227.050 0.835 2232.190 4.280 ;
        RECT 2233.030 0.835 2238.170 4.280 ;
        RECT 2239.010 0.835 2244.150 4.280 ;
        RECT 2244.990 0.835 2250.130 4.280 ;
        RECT 2250.970 0.835 2256.110 4.280 ;
        RECT 2256.950 0.835 2262.090 4.280 ;
        RECT 2262.930 0.835 2268.070 4.280 ;
        RECT 2268.910 0.835 2274.050 4.280 ;
        RECT 2274.890 0.835 2280.030 4.280 ;
        RECT 2280.870 0.835 2286.010 4.280 ;
        RECT 2286.850 0.835 2291.990 4.280 ;
        RECT 2292.830 0.835 2297.970 4.280 ;
        RECT 2298.810 0.835 2303.950 4.280 ;
        RECT 2304.790 0.835 2309.930 4.280 ;
        RECT 2310.770 0.835 2315.910 4.280 ;
        RECT 2316.750 0.835 2321.890 4.280 ;
        RECT 2322.730 0.835 2327.870 4.280 ;
        RECT 2328.710 0.835 2333.850 4.280 ;
        RECT 2334.690 0.835 2339.830 4.280 ;
        RECT 2340.670 0.835 2345.810 4.280 ;
        RECT 2346.650 0.835 2351.790 4.280 ;
        RECT 2352.630 0.835 2357.770 4.280 ;
        RECT 2358.610 0.835 2363.750 4.280 ;
        RECT 2364.590 0.835 2369.730 4.280 ;
        RECT 2370.570 0.835 2375.710 4.280 ;
        RECT 2376.550 0.835 2381.690 4.280 ;
        RECT 2382.530 0.835 2387.670 4.280 ;
        RECT 2388.510 0.835 2393.650 4.280 ;
        RECT 2394.490 0.835 2399.630 4.280 ;
        RECT 2400.470 0.835 2405.610 4.280 ;
        RECT 2406.450 0.835 2411.590 4.280 ;
        RECT 2412.430 0.835 2417.570 4.280 ;
        RECT 2418.410 0.835 2423.550 4.280 ;
        RECT 2424.390 0.835 2429.530 4.280 ;
        RECT 2430.370 0.835 2435.510 4.280 ;
        RECT 2436.350 0.835 2441.490 4.280 ;
        RECT 2442.330 0.835 2447.470 4.280 ;
        RECT 2448.310 0.835 2453.450 4.280 ;
        RECT 2454.290 0.835 2459.430 4.280 ;
        RECT 2460.270 0.835 2465.410 4.280 ;
        RECT 2466.250 0.835 2471.390 4.280 ;
        RECT 2472.230 0.835 2477.370 4.280 ;
        RECT 2478.210 0.835 2483.350 4.280 ;
        RECT 2484.190 0.835 2489.330 4.280 ;
        RECT 2490.170 0.835 2495.310 4.280 ;
        RECT 2496.150 0.835 2501.290 4.280 ;
        RECT 2502.130 0.835 2507.270 4.280 ;
        RECT 2508.110 0.835 2513.250 4.280 ;
        RECT 2514.090 0.835 2519.230 4.280 ;
        RECT 2520.070 0.835 2525.210 4.280 ;
        RECT 2526.050 0.835 2531.190 4.280 ;
        RECT 2532.030 0.835 2537.170 4.280 ;
        RECT 2538.010 0.835 2543.150 4.280 ;
        RECT 2543.990 0.835 2549.130 4.280 ;
        RECT 2549.970 0.835 2555.110 4.280 ;
        RECT 2555.950 0.835 2561.090 4.280 ;
        RECT 2561.930 0.835 2567.070 4.280 ;
        RECT 2567.910 0.835 2573.050 4.280 ;
        RECT 2573.890 0.835 2579.030 4.280 ;
        RECT 2579.870 0.835 2585.010 4.280 ;
        RECT 2585.850 0.835 2590.990 4.280 ;
        RECT 2591.830 0.835 2596.970 4.280 ;
        RECT 2597.810 0.835 2602.950 4.280 ;
        RECT 2603.790 0.835 2608.930 4.280 ;
        RECT 2609.770 0.835 2614.910 4.280 ;
        RECT 2615.750 0.835 2620.890 4.280 ;
        RECT 2621.730 0.835 2626.870 4.280 ;
        RECT 2627.710 0.835 2632.850 4.280 ;
        RECT 2633.690 0.835 2638.830 4.280 ;
        RECT 2639.670 0.835 2644.810 4.280 ;
        RECT 2645.650 0.835 2650.790 4.280 ;
        RECT 2651.630 0.835 2656.770 4.280 ;
        RECT 2657.610 0.835 2662.750 4.280 ;
        RECT 2663.590 0.835 2668.730 4.280 ;
        RECT 2669.570 0.835 2674.710 4.280 ;
        RECT 2675.550 0.835 2680.690 4.280 ;
        RECT 2681.530 0.835 2686.670 4.280 ;
        RECT 2687.510 0.835 2692.650 4.280 ;
        RECT 2693.490 0.835 2698.630 4.280 ;
        RECT 2699.470 0.835 2704.610 4.280 ;
        RECT 2705.450 0.835 2710.590 4.280 ;
        RECT 2711.430 0.835 2716.570 4.280 ;
        RECT 2717.410 0.835 2722.550 4.280 ;
        RECT 2723.390 0.835 2728.530 4.280 ;
        RECT 2729.370 0.835 2734.510 4.280 ;
        RECT 2735.350 0.835 2740.490 4.280 ;
        RECT 2741.330 0.835 2746.470 4.280 ;
        RECT 2747.310 0.835 2752.450 4.280 ;
        RECT 2753.290 0.835 2758.430 4.280 ;
        RECT 2759.270 0.835 2764.410 4.280 ;
        RECT 2765.250 0.835 2770.390 4.280 ;
        RECT 2771.230 0.835 2776.370 4.280 ;
        RECT 2777.210 0.835 2782.350 4.280 ;
        RECT 2783.190 0.835 2788.330 4.280 ;
        RECT 2789.170 0.835 2794.310 4.280 ;
        RECT 2795.150 0.835 2800.290 4.280 ;
        RECT 2801.130 0.835 2806.270 4.280 ;
        RECT 2807.110 0.835 2812.250 4.280 ;
        RECT 2813.090 0.835 2818.230 4.280 ;
        RECT 2819.070 0.835 2824.210 4.280 ;
        RECT 2825.050 0.835 2830.190 4.280 ;
        RECT 2831.030 0.835 2836.170 4.280 ;
        RECT 2837.010 0.835 2842.150 4.280 ;
        RECT 2842.990 0.835 2848.130 4.280 ;
        RECT 2848.970 0.835 2854.110 4.280 ;
        RECT 2854.950 0.835 2860.090 4.280 ;
        RECT 2860.930 0.835 2866.070 4.280 ;
        RECT 2866.910 0.835 2872.050 4.280 ;
        RECT 2872.890 0.835 2878.030 4.280 ;
        RECT 2878.870 0.835 2884.010 4.280 ;
        RECT 2884.850 0.835 2889.990 4.280 ;
        RECT 2890.830 0.835 2895.970 4.280 ;
        RECT 2896.810 0.835 2901.950 4.280 ;
        RECT 2902.790 0.835 2907.930 4.280 ;
        RECT 2908.770 0.835 2913.910 4.280 ;
        RECT 2914.750 0.835 2919.890 4.280 ;
        RECT 2920.730 0.835 2925.870 4.280 ;
        RECT 2926.710 0.835 2931.850 4.280 ;
        RECT 2932.690 0.835 2937.830 4.280 ;
        RECT 2938.670 0.835 2943.810 4.280 ;
        RECT 2944.650 0.835 2949.790 4.280 ;
        RECT 2950.630 0.835 2955.770 4.280 ;
        RECT 2956.610 0.835 2961.750 4.280 ;
        RECT 2962.590 0.835 2967.730 4.280 ;
        RECT 2968.570 0.835 2973.710 4.280 ;
        RECT 2974.550 0.835 2997.730 4.280 ;
      LAYER met3 ;
        RECT 4.000 3548.600 3002.000 3585.125 ;
        RECT 4.000 3547.200 3001.600 3548.600 ;
        RECT 4.000 3541.120 3002.000 3547.200 ;
        RECT 4.400 3539.720 3002.000 3541.120 ;
        RECT 4.000 3469.040 3002.000 3539.720 ;
        RECT 4.000 3467.640 3001.600 3469.040 ;
        RECT 4.000 3456.120 3002.000 3467.640 ;
        RECT 4.400 3454.720 3002.000 3456.120 ;
        RECT 4.000 3389.480 3002.000 3454.720 ;
        RECT 4.000 3388.080 3001.600 3389.480 ;
        RECT 4.000 3371.120 3002.000 3388.080 ;
        RECT 4.400 3369.720 3002.000 3371.120 ;
        RECT 4.000 3309.920 3002.000 3369.720 ;
        RECT 4.000 3308.520 3001.600 3309.920 ;
        RECT 4.000 3286.120 3002.000 3308.520 ;
        RECT 4.400 3284.720 3002.000 3286.120 ;
        RECT 4.000 3230.360 3002.000 3284.720 ;
        RECT 4.000 3228.960 3001.600 3230.360 ;
        RECT 4.000 3201.120 3002.000 3228.960 ;
        RECT 4.400 3199.720 3002.000 3201.120 ;
        RECT 4.000 3150.800 3002.000 3199.720 ;
        RECT 4.000 3149.400 3001.600 3150.800 ;
        RECT 4.000 3116.120 3002.000 3149.400 ;
        RECT 4.400 3114.720 3002.000 3116.120 ;
        RECT 4.000 3071.240 3002.000 3114.720 ;
        RECT 4.000 3069.840 3001.600 3071.240 ;
        RECT 4.000 3031.120 3002.000 3069.840 ;
        RECT 4.400 3029.720 3002.000 3031.120 ;
        RECT 4.000 2991.680 3002.000 3029.720 ;
        RECT 4.000 2990.280 3001.600 2991.680 ;
        RECT 4.000 2946.120 3002.000 2990.280 ;
        RECT 4.400 2944.720 3002.000 2946.120 ;
        RECT 4.000 2912.120 3002.000 2944.720 ;
        RECT 4.000 2910.720 3001.600 2912.120 ;
        RECT 4.000 2861.120 3002.000 2910.720 ;
        RECT 4.400 2859.720 3002.000 2861.120 ;
        RECT 4.000 2832.560 3002.000 2859.720 ;
        RECT 4.000 2831.160 3001.600 2832.560 ;
        RECT 4.000 2776.120 3002.000 2831.160 ;
        RECT 4.400 2774.720 3002.000 2776.120 ;
        RECT 4.000 2753.000 3002.000 2774.720 ;
        RECT 4.000 2751.600 3001.600 2753.000 ;
        RECT 4.000 2691.120 3002.000 2751.600 ;
        RECT 4.400 2689.720 3002.000 2691.120 ;
        RECT 4.000 2673.440 3002.000 2689.720 ;
        RECT 4.000 2672.040 3001.600 2673.440 ;
        RECT 4.000 2606.120 3002.000 2672.040 ;
        RECT 4.400 2604.720 3002.000 2606.120 ;
        RECT 4.000 2593.880 3002.000 2604.720 ;
        RECT 4.000 2592.480 3001.600 2593.880 ;
        RECT 4.000 2521.120 3002.000 2592.480 ;
        RECT 4.400 2519.720 3002.000 2521.120 ;
        RECT 4.000 2514.320 3002.000 2519.720 ;
        RECT 4.000 2512.920 3001.600 2514.320 ;
        RECT 4.000 2436.120 3002.000 2512.920 ;
        RECT 4.400 2434.760 3002.000 2436.120 ;
        RECT 4.400 2434.720 3001.600 2434.760 ;
        RECT 4.000 2433.360 3001.600 2434.720 ;
        RECT 4.000 2355.200 3002.000 2433.360 ;
        RECT 4.000 2353.800 3001.600 2355.200 ;
        RECT 4.000 2351.120 3002.000 2353.800 ;
        RECT 4.400 2349.720 3002.000 2351.120 ;
        RECT 4.000 2275.640 3002.000 2349.720 ;
        RECT 4.000 2274.240 3001.600 2275.640 ;
        RECT 4.000 2266.120 3002.000 2274.240 ;
        RECT 4.400 2264.720 3002.000 2266.120 ;
        RECT 4.000 2196.080 3002.000 2264.720 ;
        RECT 4.000 2194.680 3001.600 2196.080 ;
        RECT 4.000 2181.120 3002.000 2194.680 ;
        RECT 4.400 2179.720 3002.000 2181.120 ;
        RECT 4.000 2116.520 3002.000 2179.720 ;
        RECT 4.000 2115.120 3001.600 2116.520 ;
        RECT 4.000 2096.120 3002.000 2115.120 ;
        RECT 4.400 2094.720 3002.000 2096.120 ;
        RECT 4.000 2036.960 3002.000 2094.720 ;
        RECT 4.000 2035.560 3001.600 2036.960 ;
        RECT 4.000 2011.120 3002.000 2035.560 ;
        RECT 4.400 2009.720 3002.000 2011.120 ;
        RECT 4.000 1957.400 3002.000 2009.720 ;
        RECT 4.000 1956.000 3001.600 1957.400 ;
        RECT 4.000 1926.120 3002.000 1956.000 ;
        RECT 4.400 1924.720 3002.000 1926.120 ;
        RECT 4.000 1877.840 3002.000 1924.720 ;
        RECT 4.000 1876.440 3001.600 1877.840 ;
        RECT 4.000 1841.120 3002.000 1876.440 ;
        RECT 4.400 1839.720 3002.000 1841.120 ;
        RECT 4.000 1798.280 3002.000 1839.720 ;
        RECT 4.000 1796.880 3001.600 1798.280 ;
        RECT 4.000 1756.120 3002.000 1796.880 ;
        RECT 4.400 1754.720 3002.000 1756.120 ;
        RECT 4.000 1718.720 3002.000 1754.720 ;
        RECT 4.000 1717.320 3001.600 1718.720 ;
        RECT 4.000 1671.120 3002.000 1717.320 ;
        RECT 4.400 1669.720 3002.000 1671.120 ;
        RECT 4.000 1639.160 3002.000 1669.720 ;
        RECT 4.000 1637.760 3001.600 1639.160 ;
        RECT 4.000 1586.120 3002.000 1637.760 ;
        RECT 4.400 1584.720 3002.000 1586.120 ;
        RECT 4.000 1559.600 3002.000 1584.720 ;
        RECT 4.000 1558.200 3001.600 1559.600 ;
        RECT 4.000 1501.120 3002.000 1558.200 ;
        RECT 4.400 1499.720 3002.000 1501.120 ;
        RECT 4.000 1480.040 3002.000 1499.720 ;
        RECT 4.000 1478.640 3001.600 1480.040 ;
        RECT 4.000 1416.120 3002.000 1478.640 ;
        RECT 4.400 1414.720 3002.000 1416.120 ;
        RECT 4.000 1400.480 3002.000 1414.720 ;
        RECT 4.000 1399.080 3001.600 1400.480 ;
        RECT 4.000 1331.120 3002.000 1399.080 ;
        RECT 4.400 1329.720 3002.000 1331.120 ;
        RECT 4.000 1320.920 3002.000 1329.720 ;
        RECT 4.000 1319.520 3001.600 1320.920 ;
        RECT 4.000 1246.120 3002.000 1319.520 ;
        RECT 4.400 1244.720 3002.000 1246.120 ;
        RECT 4.000 1241.360 3002.000 1244.720 ;
        RECT 4.000 1239.960 3001.600 1241.360 ;
        RECT 4.000 1161.800 3002.000 1239.960 ;
        RECT 4.000 1161.120 3001.600 1161.800 ;
        RECT 4.400 1160.400 3001.600 1161.120 ;
        RECT 4.400 1159.720 3002.000 1160.400 ;
        RECT 4.000 1082.240 3002.000 1159.720 ;
        RECT 4.000 1080.840 3001.600 1082.240 ;
        RECT 4.000 1076.120 3002.000 1080.840 ;
        RECT 4.400 1074.720 3002.000 1076.120 ;
        RECT 4.000 1002.680 3002.000 1074.720 ;
        RECT 4.000 1001.280 3001.600 1002.680 ;
        RECT 4.000 991.120 3002.000 1001.280 ;
        RECT 4.400 989.720 3002.000 991.120 ;
        RECT 4.000 923.120 3002.000 989.720 ;
        RECT 4.000 921.720 3001.600 923.120 ;
        RECT 4.000 906.120 3002.000 921.720 ;
        RECT 4.400 904.720 3002.000 906.120 ;
        RECT 4.000 843.560 3002.000 904.720 ;
        RECT 4.000 842.160 3001.600 843.560 ;
        RECT 4.000 821.120 3002.000 842.160 ;
        RECT 4.400 819.720 3002.000 821.120 ;
        RECT 4.000 764.000 3002.000 819.720 ;
        RECT 4.000 762.600 3001.600 764.000 ;
        RECT 4.000 736.120 3002.000 762.600 ;
        RECT 4.400 734.720 3002.000 736.120 ;
        RECT 4.000 684.440 3002.000 734.720 ;
        RECT 4.000 683.040 3001.600 684.440 ;
        RECT 4.000 651.120 3002.000 683.040 ;
        RECT 4.400 649.720 3002.000 651.120 ;
        RECT 4.000 604.880 3002.000 649.720 ;
        RECT 4.000 603.480 3001.600 604.880 ;
        RECT 4.000 566.120 3002.000 603.480 ;
        RECT 4.400 564.720 3002.000 566.120 ;
        RECT 4.000 525.320 3002.000 564.720 ;
        RECT 4.000 523.920 3001.600 525.320 ;
        RECT 4.000 481.120 3002.000 523.920 ;
        RECT 4.400 479.720 3002.000 481.120 ;
        RECT 4.000 445.760 3002.000 479.720 ;
        RECT 4.000 444.360 3001.600 445.760 ;
        RECT 4.000 396.120 3002.000 444.360 ;
        RECT 4.400 394.720 3002.000 396.120 ;
        RECT 4.000 366.200 3002.000 394.720 ;
        RECT 4.000 364.800 3001.600 366.200 ;
        RECT 4.000 311.120 3002.000 364.800 ;
        RECT 4.400 309.720 3002.000 311.120 ;
        RECT 4.000 286.640 3002.000 309.720 ;
        RECT 4.000 285.240 3001.600 286.640 ;
        RECT 4.000 226.120 3002.000 285.240 ;
        RECT 4.400 224.720 3002.000 226.120 ;
        RECT 4.000 207.080 3002.000 224.720 ;
        RECT 4.000 205.680 3001.600 207.080 ;
        RECT 4.000 141.120 3002.000 205.680 ;
        RECT 4.400 139.720 3002.000 141.120 ;
        RECT 4.000 127.520 3002.000 139.720 ;
        RECT 4.000 126.120 3001.600 127.520 ;
        RECT 4.000 56.120 3002.000 126.120 ;
        RECT 4.400 54.720 3002.000 56.120 ;
        RECT 4.000 47.960 3002.000 54.720 ;
        RECT 4.000 46.560 3001.600 47.960 ;
        RECT 4.000 0.855 3002.000 46.560 ;
      LAYER met4 ;
        RECT 10.910 2.895 12.440 3583.425 ;
        RECT 31.240 3531.200 89.240 3583.425 ;
        RECT 31.240 2904.320 37.980 3531.200 ;
        RECT 56.780 3525.600 89.240 3531.200 ;
        RECT 108.040 3525.600 166.040 3583.425 ;
        RECT 184.840 3525.600 242.840 3583.425 ;
        RECT 261.640 3525.600 319.640 3583.425 ;
        RECT 338.440 3525.600 396.440 3583.425 ;
        RECT 415.240 3525.600 473.240 3583.425 ;
        RECT 492.040 3525.600 550.040 3583.425 ;
        RECT 568.840 3525.600 626.840 3583.425 ;
        RECT 645.640 3525.600 703.640 3583.425 ;
        RECT 722.440 3525.600 780.440 3583.425 ;
        RECT 799.240 3525.600 857.240 3583.425 ;
        RECT 876.040 3525.600 934.040 3583.425 ;
        RECT 952.840 3525.600 1010.840 3583.425 ;
        RECT 1029.640 3528.480 1087.640 3583.425 ;
        RECT 56.780 2906.400 1010.840 3525.600 ;
        RECT 56.780 2904.320 89.240 2906.400 ;
        RECT 31.240 2829.440 89.240 2904.320 ;
        RECT 31.240 2202.560 37.980 2829.440 ;
        RECT 56.780 2826.600 89.240 2829.440 ;
        RECT 108.040 2826.600 166.040 2906.400 ;
        RECT 184.840 2826.600 242.840 2906.400 ;
        RECT 261.640 2826.600 319.640 2906.400 ;
        RECT 338.440 2826.600 396.440 2906.400 ;
        RECT 415.240 2826.600 473.240 2906.400 ;
        RECT 492.040 2826.600 550.040 2906.400 ;
        RECT 568.840 2826.600 626.840 2906.400 ;
        RECT 645.640 2826.600 703.640 2906.400 ;
        RECT 722.440 2826.600 780.440 2906.400 ;
        RECT 799.240 2826.600 857.240 2906.400 ;
        RECT 876.040 2826.600 934.040 2906.400 ;
        RECT 952.840 2826.600 1010.840 2906.400 ;
        RECT 1039.440 3525.600 1087.640 3528.480 ;
        RECT 1106.440 3525.600 1164.440 3583.425 ;
        RECT 1183.240 3525.600 1241.240 3583.425 ;
        RECT 1260.040 3525.600 1318.040 3583.425 ;
        RECT 1336.840 3525.600 1394.840 3583.425 ;
        RECT 1413.640 3525.600 1471.640 3583.425 ;
        RECT 1490.440 3525.600 1548.440 3583.425 ;
        RECT 1567.240 3525.600 1625.240 3583.425 ;
        RECT 1644.040 3525.600 1702.040 3583.425 ;
        RECT 1720.840 3525.600 1778.840 3583.425 ;
        RECT 1797.640 3525.600 1855.640 3583.425 ;
        RECT 1874.440 3525.600 1932.440 3583.425 ;
        RECT 1951.240 3531.200 2009.240 3583.425 ;
        RECT 1951.240 3525.600 1969.880 3531.200 ;
        RECT 1039.440 2906.400 1969.880 3525.600 ;
        RECT 1039.440 2901.600 1087.640 2906.400 ;
        RECT 1029.640 2846.200 1087.640 2901.600 ;
        RECT 56.780 2207.400 1010.840 2826.600 ;
        RECT 56.780 2202.560 89.240 2207.400 ;
        RECT 31.240 2133.120 89.240 2202.560 ;
        RECT 31.240 1506.240 37.980 2133.120 ;
        RECT 56.780 2127.600 89.240 2133.120 ;
        RECT 108.040 2127.600 166.040 2207.400 ;
        RECT 184.840 2127.600 242.840 2207.400 ;
        RECT 261.640 2127.600 319.640 2207.400 ;
        RECT 338.440 2127.600 396.440 2207.400 ;
        RECT 415.240 2127.600 473.240 2207.400 ;
        RECT 492.040 2127.600 550.040 2207.400 ;
        RECT 568.840 2127.600 626.840 2207.400 ;
        RECT 645.640 2127.600 703.640 2207.400 ;
        RECT 722.440 2127.600 780.440 2207.400 ;
        RECT 799.240 2127.600 857.240 2207.400 ;
        RECT 876.040 2127.600 934.040 2207.400 ;
        RECT 952.840 2127.600 1010.840 2207.400 ;
        RECT 1039.440 2826.600 1087.640 2846.200 ;
        RECT 1106.440 2826.600 1164.440 2906.400 ;
        RECT 1183.240 2826.600 1241.240 2906.400 ;
        RECT 1260.040 2826.600 1318.040 2906.400 ;
        RECT 1336.840 2826.600 1394.840 2906.400 ;
        RECT 1413.640 2826.600 1471.640 2906.400 ;
        RECT 1490.440 2826.600 1548.440 2906.400 ;
        RECT 1567.240 2826.600 1625.240 2906.400 ;
        RECT 1644.040 2826.600 1702.040 2906.400 ;
        RECT 1720.840 2826.600 1778.840 2906.400 ;
        RECT 1797.640 2826.600 1855.640 2906.400 ;
        RECT 1874.440 2826.600 1932.440 2906.400 ;
        RECT 1951.240 2901.600 1969.880 2906.400 ;
        RECT 1979.680 2901.600 1980.000 3531.200 ;
        RECT 1989.800 3525.600 2009.240 3531.200 ;
        RECT 2028.040 3525.600 2086.040 3583.425 ;
        RECT 2104.840 3525.600 2162.840 3583.425 ;
        RECT 2181.640 3525.600 2239.640 3583.425 ;
        RECT 2258.440 3525.600 2316.440 3583.425 ;
        RECT 2335.240 3525.600 2393.240 3583.425 ;
        RECT 2412.040 3525.600 2470.040 3583.425 ;
        RECT 2488.840 3525.600 2546.840 3583.425 ;
        RECT 2565.640 3525.600 2623.640 3583.425 ;
        RECT 2642.440 3525.600 2700.440 3583.425 ;
        RECT 2719.240 3525.600 2777.240 3583.425 ;
        RECT 2796.040 3525.600 2854.040 3583.425 ;
        RECT 2872.840 3525.600 2930.840 3583.425 ;
        RECT 1989.800 2906.400 2930.840 3525.600 ;
        RECT 1989.800 2901.600 2009.240 2906.400 ;
        RECT 1951.240 2846.200 2009.240 2901.600 ;
        RECT 1951.240 2826.600 1969.880 2846.200 ;
        RECT 1039.440 2207.400 1969.880 2826.600 ;
        RECT 1039.440 2205.280 1087.640 2207.400 ;
        RECT 1029.640 2130.400 1087.640 2205.280 ;
        RECT 56.780 1508.400 1010.840 2127.600 ;
        RECT 56.780 1506.240 89.240 1508.400 ;
        RECT 31.240 1431.360 89.240 1506.240 ;
        RECT 31.240 804.480 37.980 1431.360 ;
        RECT 56.780 1428.600 89.240 1431.360 ;
        RECT 108.040 1428.600 166.040 1508.400 ;
        RECT 184.840 1428.600 242.840 1508.400 ;
        RECT 261.640 1428.600 319.640 1508.400 ;
        RECT 338.440 1428.600 396.440 1508.400 ;
        RECT 415.240 1428.600 473.240 1508.400 ;
        RECT 492.040 1428.600 550.040 1508.400 ;
        RECT 568.840 1428.600 626.840 1508.400 ;
        RECT 645.640 1428.600 703.640 1508.400 ;
        RECT 722.440 1428.600 780.440 1508.400 ;
        RECT 799.240 1428.600 857.240 1508.400 ;
        RECT 876.040 1428.600 934.040 1508.400 ;
        RECT 952.840 1428.600 1010.840 1508.400 ;
        RECT 1039.440 2127.600 1087.640 2130.400 ;
        RECT 1106.440 2127.600 1164.440 2207.400 ;
        RECT 1183.240 2127.600 1241.240 2207.400 ;
        RECT 1260.040 2127.600 1318.040 2207.400 ;
        RECT 1336.840 2127.600 1394.840 2207.400 ;
        RECT 1413.640 2127.600 1471.640 2207.400 ;
        RECT 1490.440 2127.600 1548.440 2207.400 ;
        RECT 1567.240 2127.600 1625.240 2207.400 ;
        RECT 1644.040 2127.600 1702.040 2207.400 ;
        RECT 1720.840 2127.600 1778.840 2207.400 ;
        RECT 1797.640 2127.600 1855.640 2207.400 ;
        RECT 1874.440 2127.600 1932.440 2207.400 ;
        RECT 1951.240 2202.560 1969.880 2207.400 ;
        RECT 1979.680 2832.160 2009.240 2846.200 ;
        RECT 1979.680 2202.560 1980.000 2832.160 ;
        RECT 1989.800 2826.600 2009.240 2832.160 ;
        RECT 2028.040 2826.600 2086.040 2906.400 ;
        RECT 2104.840 2826.600 2162.840 2906.400 ;
        RECT 2181.640 2826.600 2239.640 2906.400 ;
        RECT 2258.440 2826.600 2316.440 2906.400 ;
        RECT 2335.240 2826.600 2393.240 2906.400 ;
        RECT 2412.040 2826.600 2470.040 2906.400 ;
        RECT 2488.840 2826.600 2546.840 2906.400 ;
        RECT 2565.640 2826.600 2623.640 2906.400 ;
        RECT 2642.440 2826.600 2700.440 2906.400 ;
        RECT 2719.240 2826.600 2777.240 2906.400 ;
        RECT 2796.040 2826.600 2854.040 2906.400 ;
        RECT 2872.840 2826.600 2930.840 2906.400 ;
        RECT 1989.800 2207.400 2930.840 2826.600 ;
        RECT 1989.800 2202.560 2009.240 2207.400 ;
        RECT 1951.240 2133.120 2009.240 2202.560 ;
        RECT 1951.240 2127.600 1969.880 2133.120 ;
        RECT 1039.440 1508.400 1969.880 2127.600 ;
        RECT 1039.440 1503.520 1087.640 1508.400 ;
        RECT 1029.640 1434.080 1087.640 1503.520 ;
        RECT 56.780 809.400 1010.840 1428.600 ;
        RECT 56.780 804.480 89.240 809.400 ;
        RECT 31.240 735.040 89.240 804.480 ;
        RECT 31.240 95.220 37.980 735.040 ;
        RECT 56.780 729.600 89.240 735.040 ;
        RECT 108.040 729.600 166.040 809.400 ;
        RECT 184.840 729.600 242.840 809.400 ;
        RECT 261.640 729.600 319.640 809.400 ;
        RECT 338.440 729.600 396.440 809.400 ;
        RECT 415.240 729.600 473.240 809.400 ;
        RECT 492.040 729.600 550.040 809.400 ;
        RECT 568.840 729.600 626.840 809.400 ;
        RECT 645.640 729.600 703.640 809.400 ;
        RECT 722.440 729.600 780.440 809.400 ;
        RECT 799.240 729.600 857.240 809.400 ;
        RECT 876.040 729.600 934.040 809.400 ;
        RECT 952.840 729.600 1010.840 809.400 ;
        RECT 1039.440 1428.600 1087.640 1434.080 ;
        RECT 1106.440 1428.600 1164.440 1508.400 ;
        RECT 1183.240 1428.600 1241.240 1508.400 ;
        RECT 1260.040 1428.600 1318.040 1508.400 ;
        RECT 1336.840 1428.600 1394.840 1508.400 ;
        RECT 1413.640 1428.600 1471.640 1508.400 ;
        RECT 1490.440 1428.600 1548.440 1508.400 ;
        RECT 1567.240 1428.600 1625.240 1508.400 ;
        RECT 1644.040 1428.600 1702.040 1508.400 ;
        RECT 1720.840 1428.600 1778.840 1508.400 ;
        RECT 1797.640 1428.600 1855.640 1508.400 ;
        RECT 1874.440 1428.600 1932.440 1508.400 ;
        RECT 1951.240 1503.520 1969.880 1508.400 ;
        RECT 1979.680 1503.520 1980.000 2133.120 ;
        RECT 1989.800 2127.600 2009.240 2133.120 ;
        RECT 2028.040 2127.600 2086.040 2207.400 ;
        RECT 2104.840 2127.600 2162.840 2207.400 ;
        RECT 2181.640 2127.600 2239.640 2207.400 ;
        RECT 2258.440 2127.600 2316.440 2207.400 ;
        RECT 2335.240 2127.600 2393.240 2207.400 ;
        RECT 2412.040 2127.600 2470.040 2207.400 ;
        RECT 2488.840 2127.600 2546.840 2207.400 ;
        RECT 2565.640 2127.600 2623.640 2207.400 ;
        RECT 2642.440 2127.600 2700.440 2207.400 ;
        RECT 2719.240 2127.600 2777.240 2207.400 ;
        RECT 2796.040 2127.600 2854.040 2207.400 ;
        RECT 2872.840 2127.600 2930.840 2207.400 ;
        RECT 1989.800 1508.400 2930.840 2127.600 ;
        RECT 1989.800 1503.520 2009.240 1508.400 ;
        RECT 1951.240 1434.080 2009.240 1503.520 ;
        RECT 1951.240 1428.600 1969.880 1434.080 ;
        RECT 1039.440 809.400 1969.880 1428.600 ;
        RECT 1039.440 807.200 1087.640 809.400 ;
        RECT 1029.640 732.320 1087.640 807.200 ;
        RECT 56.780 110.400 1010.840 729.600 ;
        RECT 56.780 95.220 89.240 110.400 ;
        RECT 31.240 2.895 89.240 95.220 ;
        RECT 108.040 2.895 166.040 110.400 ;
        RECT 184.840 2.895 242.840 110.400 ;
        RECT 261.640 2.895 319.640 110.400 ;
        RECT 338.440 2.895 396.440 110.400 ;
        RECT 415.240 2.895 473.240 110.400 ;
        RECT 492.040 2.895 550.040 110.400 ;
        RECT 568.840 2.895 626.840 110.400 ;
        RECT 645.640 2.895 703.640 110.400 ;
        RECT 722.440 2.895 780.440 110.400 ;
        RECT 799.240 2.895 857.240 110.400 ;
        RECT 876.040 2.895 934.040 110.400 ;
        RECT 952.840 2.895 1010.840 110.400 ;
        RECT 1039.440 729.600 1087.640 732.320 ;
        RECT 1106.440 729.600 1164.440 809.400 ;
        RECT 1183.240 729.600 1241.240 809.400 ;
        RECT 1260.040 729.600 1318.040 809.400 ;
        RECT 1336.840 729.600 1394.840 809.400 ;
        RECT 1413.640 729.600 1471.640 809.400 ;
        RECT 1490.440 729.600 1548.440 809.400 ;
        RECT 1567.240 729.600 1625.240 809.400 ;
        RECT 1644.040 729.600 1702.040 809.400 ;
        RECT 1720.840 729.600 1778.840 809.400 ;
        RECT 1797.640 729.600 1855.640 809.400 ;
        RECT 1874.440 729.600 1932.440 809.400 ;
        RECT 1951.240 804.480 1969.880 809.400 ;
        RECT 1979.680 804.480 1980.000 1434.080 ;
        RECT 1989.800 1428.600 2009.240 1434.080 ;
        RECT 2028.040 1428.600 2086.040 1508.400 ;
        RECT 2104.840 1428.600 2162.840 1508.400 ;
        RECT 2181.640 1428.600 2239.640 1508.400 ;
        RECT 2258.440 1428.600 2316.440 1508.400 ;
        RECT 2335.240 1428.600 2393.240 1508.400 ;
        RECT 2412.040 1428.600 2470.040 1508.400 ;
        RECT 2488.840 1428.600 2546.840 1508.400 ;
        RECT 2565.640 1428.600 2623.640 1508.400 ;
        RECT 2642.440 1428.600 2700.440 1508.400 ;
        RECT 2719.240 1428.600 2777.240 1508.400 ;
        RECT 2796.040 1428.600 2854.040 1508.400 ;
        RECT 2872.840 1428.600 2930.840 1508.400 ;
        RECT 1989.800 809.400 2930.840 1428.600 ;
        RECT 1989.800 804.480 2009.240 809.400 ;
        RECT 1951.240 735.040 2009.240 804.480 ;
        RECT 1951.240 729.600 1969.880 735.040 ;
        RECT 1039.440 110.400 1969.880 729.600 ;
        RECT 1039.440 105.440 1087.640 110.400 ;
        RECT 1029.640 2.895 1087.640 105.440 ;
        RECT 1106.440 2.895 1164.440 110.400 ;
        RECT 1183.240 2.895 1241.240 110.400 ;
        RECT 1260.040 2.895 1318.040 110.400 ;
        RECT 1336.840 2.895 1394.840 110.400 ;
        RECT 1413.640 2.895 1471.640 110.400 ;
        RECT 1490.440 2.895 1548.440 110.400 ;
        RECT 1567.240 2.895 1625.240 110.400 ;
        RECT 1644.040 2.895 1702.040 110.400 ;
        RECT 1720.840 2.895 1778.840 110.400 ;
        RECT 1797.640 2.895 1855.640 110.400 ;
        RECT 1874.440 2.895 1932.440 110.400 ;
        RECT 1951.240 105.440 1969.880 110.400 ;
        RECT 1979.680 105.440 1980.000 735.040 ;
        RECT 1951.240 95.220 1980.000 105.440 ;
        RECT 1989.800 729.600 2009.240 735.040 ;
        RECT 2028.040 729.600 2086.040 809.400 ;
        RECT 2104.840 729.600 2162.840 809.400 ;
        RECT 2181.640 729.600 2239.640 809.400 ;
        RECT 2258.440 729.600 2316.440 809.400 ;
        RECT 2335.240 729.600 2393.240 809.400 ;
        RECT 2412.040 729.600 2470.040 809.400 ;
        RECT 2488.840 729.600 2546.840 809.400 ;
        RECT 2565.640 729.600 2623.640 809.400 ;
        RECT 2642.440 729.600 2700.440 809.400 ;
        RECT 2719.240 729.600 2777.240 809.400 ;
        RECT 2796.040 729.600 2854.040 809.400 ;
        RECT 2872.840 729.600 2930.840 809.400 ;
        RECT 1989.800 110.400 2930.840 729.600 ;
        RECT 1989.800 95.220 2009.240 110.400 ;
        RECT 1951.240 2.895 2009.240 95.220 ;
        RECT 2028.040 2.895 2086.040 110.400 ;
        RECT 2104.840 2.895 2162.840 110.400 ;
        RECT 2181.640 2.895 2239.640 110.400 ;
        RECT 2258.440 2.895 2316.440 110.400 ;
        RECT 2335.240 2.895 2393.240 110.400 ;
        RECT 2412.040 2.895 2470.040 110.400 ;
        RECT 2488.840 2.895 2546.840 110.400 ;
        RECT 2565.640 2.895 2623.640 110.400 ;
        RECT 2642.440 2.895 2700.440 110.400 ;
        RECT 2719.240 2.895 2777.240 110.400 ;
        RECT 2796.040 2.895 2854.040 110.400 ;
        RECT 2872.840 2.895 2930.840 110.400 ;
        RECT 2949.640 3531.200 2990.130 3583.425 ;
        RECT 2949.640 2904.320 2970.020 3531.200 ;
        RECT 2988.820 2904.320 2990.130 3531.200 ;
        RECT 2949.640 2829.440 2990.130 2904.320 ;
        RECT 2949.640 2202.560 2970.020 2829.440 ;
        RECT 2988.820 2202.560 2990.130 2829.440 ;
        RECT 2949.640 2133.120 2990.130 2202.560 ;
        RECT 2949.640 1506.240 2970.020 2133.120 ;
        RECT 2988.820 1506.240 2990.130 2133.120 ;
        RECT 2949.640 1431.360 2990.130 1506.240 ;
        RECT 2949.640 804.480 2970.020 1431.360 ;
        RECT 2988.820 804.480 2990.130 1431.360 ;
        RECT 2949.640 735.040 2990.130 804.480 ;
        RECT 2949.640 95.220 2970.020 735.040 ;
        RECT 2988.820 95.220 2990.130 735.040 ;
        RECT 2949.640 2.895 2990.130 95.220 ;
      LAYER met5 ;
        RECT 10.700 3254.410 2990.340 3276.700 ;
        RECT 10.700 3177.820 2990.340 3234.210 ;
        RECT 10.700 3101.230 2990.340 3157.620 ;
        RECT 10.700 3024.640 2990.340 3081.030 ;
        RECT 10.700 2948.050 2990.340 3004.440 ;
        RECT 10.700 2871.460 2990.340 2927.850 ;
        RECT 10.700 2847.400 2990.340 2851.260 ;
        RECT 10.700 2827.200 11.240 2847.400 ;
        RECT 2950.840 2827.200 2990.340 2847.400 ;
        RECT 10.700 2794.870 2990.340 2827.200 ;
        RECT 10.700 2718.280 2990.340 2774.670 ;
        RECT 10.700 2641.690 2990.340 2698.080 ;
        RECT 10.700 2565.100 2990.340 2621.490 ;
        RECT 10.700 2488.510 2990.340 2544.900 ;
        RECT 10.700 2411.920 2990.340 2468.310 ;
        RECT 10.700 2335.330 2990.340 2391.720 ;
        RECT 10.700 2258.740 2990.340 2315.130 ;
        RECT 10.700 2182.150 2990.340 2238.540 ;
        RECT 10.700 2157.200 2990.340 2161.950 ;
        RECT 10.700 2105.560 2990.340 2137.000 ;
        RECT 10.700 2028.970 2990.340 2085.360 ;
        RECT 10.700 1952.380 2990.340 2008.770 ;
        RECT 10.700 1875.790 2990.340 1932.180 ;
        RECT 10.700 1799.200 2990.340 1855.590 ;
        RECT 10.700 1722.610 2990.340 1779.000 ;
        RECT 10.700 1646.020 2990.340 1702.410 ;
        RECT 10.700 1569.430 2990.340 1625.820 ;
        RECT 10.700 1492.840 2990.340 1549.230 ;
        RECT 10.700 1460.200 2990.340 1472.640 ;
        RECT 10.700 1440.000 11.240 1460.200 ;
        RECT 2950.840 1440.000 2990.340 1460.200 ;
        RECT 10.700 1416.250 2990.340 1440.000 ;
        RECT 10.700 1339.660 2990.340 1396.050 ;
        RECT 10.700 1263.070 2990.340 1319.460 ;
        RECT 10.700 1186.480 2990.340 1242.870 ;
        RECT 10.700 1109.890 2990.340 1166.280 ;
        RECT 10.700 1033.300 2990.340 1089.690 ;
        RECT 10.700 956.710 2990.340 1013.100 ;
        RECT 10.700 880.120 2990.340 936.510 ;
        RECT 10.700 803.530 2990.340 859.920 ;
        RECT 10.700 780.200 2990.340 783.330 ;
        RECT 10.700 726.940 2990.340 760.000 ;
        RECT 10.700 650.350 2990.340 706.740 ;
        RECT 10.700 573.760 2990.340 630.150 ;
        RECT 10.700 497.170 2990.340 553.560 ;
        RECT 10.700 420.580 2990.340 476.970 ;
        RECT 10.700 343.990 2990.340 400.380 ;
        RECT 10.700 267.400 2990.340 323.790 ;
        RECT 10.700 190.810 2990.340 247.200 ;
        RECT 10.700 114.220 2990.340 170.610 ;
        RECT 10.700 37.630 2990.340 94.020 ;
        RECT 10.700 7.700 2990.340 17.430 ;
  END
END chaos_automaton
END LIBRARY

