magic
tech sky130B
magscale 1 2
timestamp 1660177439
<< obsli1 >>
rect 1104 2159 600024 717009
<< obsm1 >>
rect 1104 280 600024 717324
<< metal2 >>
rect 11150 718400 11206 719200
rect 33414 718400 33470 719200
rect 55678 718400 55734 719200
rect 77942 718400 77998 719200
rect 100206 718400 100262 719200
rect 122470 718400 122526 719200
rect 144734 718400 144790 719200
rect 166998 718400 167054 719200
rect 189262 718400 189318 719200
rect 211526 718400 211582 719200
rect 233790 718400 233846 719200
rect 256054 718400 256110 719200
rect 278318 718400 278374 719200
rect 300582 718400 300638 719200
rect 322846 718400 322902 719200
rect 345110 718400 345166 719200
rect 367374 718400 367430 719200
rect 389638 718400 389694 719200
rect 411902 718400 411958 719200
rect 434166 718400 434222 719200
rect 456430 718400 456486 719200
rect 478694 718400 478750 719200
rect 500958 718400 501014 719200
rect 523222 718400 523278 719200
rect 545486 718400 545542 719200
rect 567750 718400 567806 719200
rect 590014 718400 590070 719200
rect 6366 0 6422 800
rect 7562 0 7618 800
rect 8758 0 8814 800
rect 9954 0 10010 800
rect 11150 0 11206 800
rect 12346 0 12402 800
rect 13542 0 13598 800
rect 14738 0 14794 800
rect 15934 0 15990 800
rect 17130 0 17186 800
rect 18326 0 18382 800
rect 19522 0 19578 800
rect 20718 0 20774 800
rect 21914 0 21970 800
rect 23110 0 23166 800
rect 24306 0 24362 800
rect 25502 0 25558 800
rect 26698 0 26754 800
rect 27894 0 27950 800
rect 29090 0 29146 800
rect 30286 0 30342 800
rect 31482 0 31538 800
rect 32678 0 32734 800
rect 33874 0 33930 800
rect 35070 0 35126 800
rect 36266 0 36322 800
rect 37462 0 37518 800
rect 38658 0 38714 800
rect 39854 0 39910 800
rect 41050 0 41106 800
rect 42246 0 42302 800
rect 43442 0 43498 800
rect 44638 0 44694 800
rect 45834 0 45890 800
rect 47030 0 47086 800
rect 48226 0 48282 800
rect 49422 0 49478 800
rect 50618 0 50674 800
rect 51814 0 51870 800
rect 53010 0 53066 800
rect 54206 0 54262 800
rect 55402 0 55458 800
rect 56598 0 56654 800
rect 57794 0 57850 800
rect 58990 0 59046 800
rect 60186 0 60242 800
rect 61382 0 61438 800
rect 62578 0 62634 800
rect 63774 0 63830 800
rect 64970 0 65026 800
rect 66166 0 66222 800
rect 67362 0 67418 800
rect 68558 0 68614 800
rect 69754 0 69810 800
rect 70950 0 71006 800
rect 72146 0 72202 800
rect 73342 0 73398 800
rect 74538 0 74594 800
rect 75734 0 75790 800
rect 76930 0 76986 800
rect 78126 0 78182 800
rect 79322 0 79378 800
rect 80518 0 80574 800
rect 81714 0 81770 800
rect 82910 0 82966 800
rect 84106 0 84162 800
rect 85302 0 85358 800
rect 86498 0 86554 800
rect 87694 0 87750 800
rect 88890 0 88946 800
rect 90086 0 90142 800
rect 91282 0 91338 800
rect 92478 0 92534 800
rect 93674 0 93730 800
rect 94870 0 94926 800
rect 96066 0 96122 800
rect 97262 0 97318 800
rect 98458 0 98514 800
rect 99654 0 99710 800
rect 100850 0 100906 800
rect 102046 0 102102 800
rect 103242 0 103298 800
rect 104438 0 104494 800
rect 105634 0 105690 800
rect 106830 0 106886 800
rect 108026 0 108082 800
rect 109222 0 109278 800
rect 110418 0 110474 800
rect 111614 0 111670 800
rect 112810 0 112866 800
rect 114006 0 114062 800
rect 115202 0 115258 800
rect 116398 0 116454 800
rect 117594 0 117650 800
rect 118790 0 118846 800
rect 119986 0 120042 800
rect 121182 0 121238 800
rect 122378 0 122434 800
rect 123574 0 123630 800
rect 124770 0 124826 800
rect 125966 0 126022 800
rect 127162 0 127218 800
rect 128358 0 128414 800
rect 129554 0 129610 800
rect 130750 0 130806 800
rect 131946 0 132002 800
rect 133142 0 133198 800
rect 134338 0 134394 800
rect 135534 0 135590 800
rect 136730 0 136786 800
rect 137926 0 137982 800
rect 139122 0 139178 800
rect 140318 0 140374 800
rect 141514 0 141570 800
rect 142710 0 142766 800
rect 143906 0 143962 800
rect 145102 0 145158 800
rect 146298 0 146354 800
rect 147494 0 147550 800
rect 148690 0 148746 800
rect 149886 0 149942 800
rect 151082 0 151138 800
rect 152278 0 152334 800
rect 153474 0 153530 800
rect 154670 0 154726 800
rect 155866 0 155922 800
rect 157062 0 157118 800
rect 158258 0 158314 800
rect 159454 0 159510 800
rect 160650 0 160706 800
rect 161846 0 161902 800
rect 163042 0 163098 800
rect 164238 0 164294 800
rect 165434 0 165490 800
rect 166630 0 166686 800
rect 167826 0 167882 800
rect 169022 0 169078 800
rect 170218 0 170274 800
rect 171414 0 171470 800
rect 172610 0 172666 800
rect 173806 0 173862 800
rect 175002 0 175058 800
rect 176198 0 176254 800
rect 177394 0 177450 800
rect 178590 0 178646 800
rect 179786 0 179842 800
rect 180982 0 181038 800
rect 182178 0 182234 800
rect 183374 0 183430 800
rect 184570 0 184626 800
rect 185766 0 185822 800
rect 186962 0 187018 800
rect 188158 0 188214 800
rect 189354 0 189410 800
rect 190550 0 190606 800
rect 191746 0 191802 800
rect 192942 0 192998 800
rect 194138 0 194194 800
rect 195334 0 195390 800
rect 196530 0 196586 800
rect 197726 0 197782 800
rect 198922 0 198978 800
rect 200118 0 200174 800
rect 201314 0 201370 800
rect 202510 0 202566 800
rect 203706 0 203762 800
rect 204902 0 204958 800
rect 206098 0 206154 800
rect 207294 0 207350 800
rect 208490 0 208546 800
rect 209686 0 209742 800
rect 210882 0 210938 800
rect 212078 0 212134 800
rect 213274 0 213330 800
rect 214470 0 214526 800
rect 215666 0 215722 800
rect 216862 0 216918 800
rect 218058 0 218114 800
rect 219254 0 219310 800
rect 220450 0 220506 800
rect 221646 0 221702 800
rect 222842 0 222898 800
rect 224038 0 224094 800
rect 225234 0 225290 800
rect 226430 0 226486 800
rect 227626 0 227682 800
rect 228822 0 228878 800
rect 230018 0 230074 800
rect 231214 0 231270 800
rect 232410 0 232466 800
rect 233606 0 233662 800
rect 234802 0 234858 800
rect 235998 0 236054 800
rect 237194 0 237250 800
rect 238390 0 238446 800
rect 239586 0 239642 800
rect 240782 0 240838 800
rect 241978 0 242034 800
rect 243174 0 243230 800
rect 244370 0 244426 800
rect 245566 0 245622 800
rect 246762 0 246818 800
rect 247958 0 248014 800
rect 249154 0 249210 800
rect 250350 0 250406 800
rect 251546 0 251602 800
rect 252742 0 252798 800
rect 253938 0 253994 800
rect 255134 0 255190 800
rect 256330 0 256386 800
rect 257526 0 257582 800
rect 258722 0 258778 800
rect 259918 0 259974 800
rect 261114 0 261170 800
rect 262310 0 262366 800
rect 263506 0 263562 800
rect 264702 0 264758 800
rect 265898 0 265954 800
rect 267094 0 267150 800
rect 268290 0 268346 800
rect 269486 0 269542 800
rect 270682 0 270738 800
rect 271878 0 271934 800
rect 273074 0 273130 800
rect 274270 0 274326 800
rect 275466 0 275522 800
rect 276662 0 276718 800
rect 277858 0 277914 800
rect 279054 0 279110 800
rect 280250 0 280306 800
rect 281446 0 281502 800
rect 282642 0 282698 800
rect 283838 0 283894 800
rect 285034 0 285090 800
rect 286230 0 286286 800
rect 287426 0 287482 800
rect 288622 0 288678 800
rect 289818 0 289874 800
rect 291014 0 291070 800
rect 292210 0 292266 800
rect 293406 0 293462 800
rect 294602 0 294658 800
rect 295798 0 295854 800
rect 296994 0 297050 800
rect 298190 0 298246 800
rect 299386 0 299442 800
rect 300582 0 300638 800
rect 301778 0 301834 800
rect 302974 0 303030 800
rect 304170 0 304226 800
rect 305366 0 305422 800
rect 306562 0 306618 800
rect 307758 0 307814 800
rect 308954 0 309010 800
rect 310150 0 310206 800
rect 311346 0 311402 800
rect 312542 0 312598 800
rect 313738 0 313794 800
rect 314934 0 314990 800
rect 316130 0 316186 800
rect 317326 0 317382 800
rect 318522 0 318578 800
rect 319718 0 319774 800
rect 320914 0 320970 800
rect 322110 0 322166 800
rect 323306 0 323362 800
rect 324502 0 324558 800
rect 325698 0 325754 800
rect 326894 0 326950 800
rect 328090 0 328146 800
rect 329286 0 329342 800
rect 330482 0 330538 800
rect 331678 0 331734 800
rect 332874 0 332930 800
rect 334070 0 334126 800
rect 335266 0 335322 800
rect 336462 0 336518 800
rect 337658 0 337714 800
rect 338854 0 338910 800
rect 340050 0 340106 800
rect 341246 0 341302 800
rect 342442 0 342498 800
rect 343638 0 343694 800
rect 344834 0 344890 800
rect 346030 0 346086 800
rect 347226 0 347282 800
rect 348422 0 348478 800
rect 349618 0 349674 800
rect 350814 0 350870 800
rect 352010 0 352066 800
rect 353206 0 353262 800
rect 354402 0 354458 800
rect 355598 0 355654 800
rect 356794 0 356850 800
rect 357990 0 358046 800
rect 359186 0 359242 800
rect 360382 0 360438 800
rect 361578 0 361634 800
rect 362774 0 362830 800
rect 363970 0 364026 800
rect 365166 0 365222 800
rect 366362 0 366418 800
rect 367558 0 367614 800
rect 368754 0 368810 800
rect 369950 0 370006 800
rect 371146 0 371202 800
rect 372342 0 372398 800
rect 373538 0 373594 800
rect 374734 0 374790 800
rect 375930 0 375986 800
rect 377126 0 377182 800
rect 378322 0 378378 800
rect 379518 0 379574 800
rect 380714 0 380770 800
rect 381910 0 381966 800
rect 383106 0 383162 800
rect 384302 0 384358 800
rect 385498 0 385554 800
rect 386694 0 386750 800
rect 387890 0 387946 800
rect 389086 0 389142 800
rect 390282 0 390338 800
rect 391478 0 391534 800
rect 392674 0 392730 800
rect 393870 0 393926 800
rect 395066 0 395122 800
rect 396262 0 396318 800
rect 397458 0 397514 800
rect 398654 0 398710 800
rect 399850 0 399906 800
rect 401046 0 401102 800
rect 402242 0 402298 800
rect 403438 0 403494 800
rect 404634 0 404690 800
rect 405830 0 405886 800
rect 407026 0 407082 800
rect 408222 0 408278 800
rect 409418 0 409474 800
rect 410614 0 410670 800
rect 411810 0 411866 800
rect 413006 0 413062 800
rect 414202 0 414258 800
rect 415398 0 415454 800
rect 416594 0 416650 800
rect 417790 0 417846 800
rect 418986 0 419042 800
rect 420182 0 420238 800
rect 421378 0 421434 800
rect 422574 0 422630 800
rect 423770 0 423826 800
rect 424966 0 425022 800
rect 426162 0 426218 800
rect 427358 0 427414 800
rect 428554 0 428610 800
rect 429750 0 429806 800
rect 430946 0 431002 800
rect 432142 0 432198 800
rect 433338 0 433394 800
rect 434534 0 434590 800
rect 435730 0 435786 800
rect 436926 0 436982 800
rect 438122 0 438178 800
rect 439318 0 439374 800
rect 440514 0 440570 800
rect 441710 0 441766 800
rect 442906 0 442962 800
rect 444102 0 444158 800
rect 445298 0 445354 800
rect 446494 0 446550 800
rect 447690 0 447746 800
rect 448886 0 448942 800
rect 450082 0 450138 800
rect 451278 0 451334 800
rect 452474 0 452530 800
rect 453670 0 453726 800
rect 454866 0 454922 800
rect 456062 0 456118 800
rect 457258 0 457314 800
rect 458454 0 458510 800
rect 459650 0 459706 800
rect 460846 0 460902 800
rect 462042 0 462098 800
rect 463238 0 463294 800
rect 464434 0 464490 800
rect 465630 0 465686 800
rect 466826 0 466882 800
rect 468022 0 468078 800
rect 469218 0 469274 800
rect 470414 0 470470 800
rect 471610 0 471666 800
rect 472806 0 472862 800
rect 474002 0 474058 800
rect 475198 0 475254 800
rect 476394 0 476450 800
rect 477590 0 477646 800
rect 478786 0 478842 800
rect 479982 0 480038 800
rect 481178 0 481234 800
rect 482374 0 482430 800
rect 483570 0 483626 800
rect 484766 0 484822 800
rect 485962 0 486018 800
rect 487158 0 487214 800
rect 488354 0 488410 800
rect 489550 0 489606 800
rect 490746 0 490802 800
rect 491942 0 491998 800
rect 493138 0 493194 800
rect 494334 0 494390 800
rect 495530 0 495586 800
rect 496726 0 496782 800
rect 497922 0 497978 800
rect 499118 0 499174 800
rect 500314 0 500370 800
rect 501510 0 501566 800
rect 502706 0 502762 800
rect 503902 0 503958 800
rect 505098 0 505154 800
rect 506294 0 506350 800
rect 507490 0 507546 800
rect 508686 0 508742 800
rect 509882 0 509938 800
rect 511078 0 511134 800
rect 512274 0 512330 800
rect 513470 0 513526 800
rect 514666 0 514722 800
rect 515862 0 515918 800
rect 517058 0 517114 800
rect 518254 0 518310 800
rect 519450 0 519506 800
rect 520646 0 520702 800
rect 521842 0 521898 800
rect 523038 0 523094 800
rect 524234 0 524290 800
rect 525430 0 525486 800
rect 526626 0 526682 800
rect 527822 0 527878 800
rect 529018 0 529074 800
rect 530214 0 530270 800
rect 531410 0 531466 800
rect 532606 0 532662 800
rect 533802 0 533858 800
rect 534998 0 535054 800
rect 536194 0 536250 800
rect 537390 0 537446 800
rect 538586 0 538642 800
rect 539782 0 539838 800
rect 540978 0 541034 800
rect 542174 0 542230 800
rect 543370 0 543426 800
rect 544566 0 544622 800
rect 545762 0 545818 800
rect 546958 0 547014 800
rect 548154 0 548210 800
rect 549350 0 549406 800
rect 550546 0 550602 800
rect 551742 0 551798 800
rect 552938 0 552994 800
rect 554134 0 554190 800
rect 555330 0 555386 800
rect 556526 0 556582 800
rect 557722 0 557778 800
rect 558918 0 558974 800
rect 560114 0 560170 800
rect 561310 0 561366 800
rect 562506 0 562562 800
rect 563702 0 563758 800
rect 564898 0 564954 800
rect 566094 0 566150 800
rect 567290 0 567346 800
rect 568486 0 568542 800
rect 569682 0 569738 800
rect 570878 0 570934 800
rect 572074 0 572130 800
rect 573270 0 573326 800
rect 574466 0 574522 800
rect 575662 0 575718 800
rect 576858 0 576914 800
rect 578054 0 578110 800
rect 579250 0 579306 800
rect 580446 0 580502 800
rect 581642 0 581698 800
rect 582838 0 582894 800
rect 584034 0 584090 800
rect 585230 0 585286 800
rect 586426 0 586482 800
rect 587622 0 587678 800
rect 588818 0 588874 800
rect 590014 0 590070 800
rect 591210 0 591266 800
rect 592406 0 592462 800
rect 593602 0 593658 800
rect 594798 0 594854 800
<< obsm2 >>
rect 1398 718344 11094 718400
rect 11262 718344 33358 718400
rect 33526 718344 55622 718400
rect 55790 718344 77886 718400
rect 78054 718344 100150 718400
rect 100318 718344 122414 718400
rect 122582 718344 144678 718400
rect 144846 718344 166942 718400
rect 167110 718344 189206 718400
rect 189374 718344 211470 718400
rect 211638 718344 233734 718400
rect 233902 718344 255998 718400
rect 256166 718344 278262 718400
rect 278430 718344 300526 718400
rect 300694 718344 322790 718400
rect 322958 718344 345054 718400
rect 345222 718344 367318 718400
rect 367486 718344 389582 718400
rect 389750 718344 411846 718400
rect 412014 718344 434110 718400
rect 434278 718344 456374 718400
rect 456542 718344 478638 718400
rect 478806 718344 500902 718400
rect 501070 718344 523166 718400
rect 523334 718344 545430 718400
rect 545598 718344 567694 718400
rect 567862 718344 589958 718400
rect 590126 718344 599546 718400
rect 1398 856 599546 718344
rect 1398 167 6310 856
rect 6478 167 7506 856
rect 7674 167 8702 856
rect 8870 167 9898 856
rect 10066 167 11094 856
rect 11262 167 12290 856
rect 12458 167 13486 856
rect 13654 167 14682 856
rect 14850 167 15878 856
rect 16046 167 17074 856
rect 17242 167 18270 856
rect 18438 167 19466 856
rect 19634 167 20662 856
rect 20830 167 21858 856
rect 22026 167 23054 856
rect 23222 167 24250 856
rect 24418 167 25446 856
rect 25614 167 26642 856
rect 26810 167 27838 856
rect 28006 167 29034 856
rect 29202 167 30230 856
rect 30398 167 31426 856
rect 31594 167 32622 856
rect 32790 167 33818 856
rect 33986 167 35014 856
rect 35182 167 36210 856
rect 36378 167 37406 856
rect 37574 167 38602 856
rect 38770 167 39798 856
rect 39966 167 40994 856
rect 41162 167 42190 856
rect 42358 167 43386 856
rect 43554 167 44582 856
rect 44750 167 45778 856
rect 45946 167 46974 856
rect 47142 167 48170 856
rect 48338 167 49366 856
rect 49534 167 50562 856
rect 50730 167 51758 856
rect 51926 167 52954 856
rect 53122 167 54150 856
rect 54318 167 55346 856
rect 55514 167 56542 856
rect 56710 167 57738 856
rect 57906 167 58934 856
rect 59102 167 60130 856
rect 60298 167 61326 856
rect 61494 167 62522 856
rect 62690 167 63718 856
rect 63886 167 64914 856
rect 65082 167 66110 856
rect 66278 167 67306 856
rect 67474 167 68502 856
rect 68670 167 69698 856
rect 69866 167 70894 856
rect 71062 167 72090 856
rect 72258 167 73286 856
rect 73454 167 74482 856
rect 74650 167 75678 856
rect 75846 167 76874 856
rect 77042 167 78070 856
rect 78238 167 79266 856
rect 79434 167 80462 856
rect 80630 167 81658 856
rect 81826 167 82854 856
rect 83022 167 84050 856
rect 84218 167 85246 856
rect 85414 167 86442 856
rect 86610 167 87638 856
rect 87806 167 88834 856
rect 89002 167 90030 856
rect 90198 167 91226 856
rect 91394 167 92422 856
rect 92590 167 93618 856
rect 93786 167 94814 856
rect 94982 167 96010 856
rect 96178 167 97206 856
rect 97374 167 98402 856
rect 98570 167 99598 856
rect 99766 167 100794 856
rect 100962 167 101990 856
rect 102158 167 103186 856
rect 103354 167 104382 856
rect 104550 167 105578 856
rect 105746 167 106774 856
rect 106942 167 107970 856
rect 108138 167 109166 856
rect 109334 167 110362 856
rect 110530 167 111558 856
rect 111726 167 112754 856
rect 112922 167 113950 856
rect 114118 167 115146 856
rect 115314 167 116342 856
rect 116510 167 117538 856
rect 117706 167 118734 856
rect 118902 167 119930 856
rect 120098 167 121126 856
rect 121294 167 122322 856
rect 122490 167 123518 856
rect 123686 167 124714 856
rect 124882 167 125910 856
rect 126078 167 127106 856
rect 127274 167 128302 856
rect 128470 167 129498 856
rect 129666 167 130694 856
rect 130862 167 131890 856
rect 132058 167 133086 856
rect 133254 167 134282 856
rect 134450 167 135478 856
rect 135646 167 136674 856
rect 136842 167 137870 856
rect 138038 167 139066 856
rect 139234 167 140262 856
rect 140430 167 141458 856
rect 141626 167 142654 856
rect 142822 167 143850 856
rect 144018 167 145046 856
rect 145214 167 146242 856
rect 146410 167 147438 856
rect 147606 167 148634 856
rect 148802 167 149830 856
rect 149998 167 151026 856
rect 151194 167 152222 856
rect 152390 167 153418 856
rect 153586 167 154614 856
rect 154782 167 155810 856
rect 155978 167 157006 856
rect 157174 167 158202 856
rect 158370 167 159398 856
rect 159566 167 160594 856
rect 160762 167 161790 856
rect 161958 167 162986 856
rect 163154 167 164182 856
rect 164350 167 165378 856
rect 165546 167 166574 856
rect 166742 167 167770 856
rect 167938 167 168966 856
rect 169134 167 170162 856
rect 170330 167 171358 856
rect 171526 167 172554 856
rect 172722 167 173750 856
rect 173918 167 174946 856
rect 175114 167 176142 856
rect 176310 167 177338 856
rect 177506 167 178534 856
rect 178702 167 179730 856
rect 179898 167 180926 856
rect 181094 167 182122 856
rect 182290 167 183318 856
rect 183486 167 184514 856
rect 184682 167 185710 856
rect 185878 167 186906 856
rect 187074 167 188102 856
rect 188270 167 189298 856
rect 189466 167 190494 856
rect 190662 167 191690 856
rect 191858 167 192886 856
rect 193054 167 194082 856
rect 194250 167 195278 856
rect 195446 167 196474 856
rect 196642 167 197670 856
rect 197838 167 198866 856
rect 199034 167 200062 856
rect 200230 167 201258 856
rect 201426 167 202454 856
rect 202622 167 203650 856
rect 203818 167 204846 856
rect 205014 167 206042 856
rect 206210 167 207238 856
rect 207406 167 208434 856
rect 208602 167 209630 856
rect 209798 167 210826 856
rect 210994 167 212022 856
rect 212190 167 213218 856
rect 213386 167 214414 856
rect 214582 167 215610 856
rect 215778 167 216806 856
rect 216974 167 218002 856
rect 218170 167 219198 856
rect 219366 167 220394 856
rect 220562 167 221590 856
rect 221758 167 222786 856
rect 222954 167 223982 856
rect 224150 167 225178 856
rect 225346 167 226374 856
rect 226542 167 227570 856
rect 227738 167 228766 856
rect 228934 167 229962 856
rect 230130 167 231158 856
rect 231326 167 232354 856
rect 232522 167 233550 856
rect 233718 167 234746 856
rect 234914 167 235942 856
rect 236110 167 237138 856
rect 237306 167 238334 856
rect 238502 167 239530 856
rect 239698 167 240726 856
rect 240894 167 241922 856
rect 242090 167 243118 856
rect 243286 167 244314 856
rect 244482 167 245510 856
rect 245678 167 246706 856
rect 246874 167 247902 856
rect 248070 167 249098 856
rect 249266 167 250294 856
rect 250462 167 251490 856
rect 251658 167 252686 856
rect 252854 167 253882 856
rect 254050 167 255078 856
rect 255246 167 256274 856
rect 256442 167 257470 856
rect 257638 167 258666 856
rect 258834 167 259862 856
rect 260030 167 261058 856
rect 261226 167 262254 856
rect 262422 167 263450 856
rect 263618 167 264646 856
rect 264814 167 265842 856
rect 266010 167 267038 856
rect 267206 167 268234 856
rect 268402 167 269430 856
rect 269598 167 270626 856
rect 270794 167 271822 856
rect 271990 167 273018 856
rect 273186 167 274214 856
rect 274382 167 275410 856
rect 275578 167 276606 856
rect 276774 167 277802 856
rect 277970 167 278998 856
rect 279166 167 280194 856
rect 280362 167 281390 856
rect 281558 167 282586 856
rect 282754 167 283782 856
rect 283950 167 284978 856
rect 285146 167 286174 856
rect 286342 167 287370 856
rect 287538 167 288566 856
rect 288734 167 289762 856
rect 289930 167 290958 856
rect 291126 167 292154 856
rect 292322 167 293350 856
rect 293518 167 294546 856
rect 294714 167 295742 856
rect 295910 167 296938 856
rect 297106 167 298134 856
rect 298302 167 299330 856
rect 299498 167 300526 856
rect 300694 167 301722 856
rect 301890 167 302918 856
rect 303086 167 304114 856
rect 304282 167 305310 856
rect 305478 167 306506 856
rect 306674 167 307702 856
rect 307870 167 308898 856
rect 309066 167 310094 856
rect 310262 167 311290 856
rect 311458 167 312486 856
rect 312654 167 313682 856
rect 313850 167 314878 856
rect 315046 167 316074 856
rect 316242 167 317270 856
rect 317438 167 318466 856
rect 318634 167 319662 856
rect 319830 167 320858 856
rect 321026 167 322054 856
rect 322222 167 323250 856
rect 323418 167 324446 856
rect 324614 167 325642 856
rect 325810 167 326838 856
rect 327006 167 328034 856
rect 328202 167 329230 856
rect 329398 167 330426 856
rect 330594 167 331622 856
rect 331790 167 332818 856
rect 332986 167 334014 856
rect 334182 167 335210 856
rect 335378 167 336406 856
rect 336574 167 337602 856
rect 337770 167 338798 856
rect 338966 167 339994 856
rect 340162 167 341190 856
rect 341358 167 342386 856
rect 342554 167 343582 856
rect 343750 167 344778 856
rect 344946 167 345974 856
rect 346142 167 347170 856
rect 347338 167 348366 856
rect 348534 167 349562 856
rect 349730 167 350758 856
rect 350926 167 351954 856
rect 352122 167 353150 856
rect 353318 167 354346 856
rect 354514 167 355542 856
rect 355710 167 356738 856
rect 356906 167 357934 856
rect 358102 167 359130 856
rect 359298 167 360326 856
rect 360494 167 361522 856
rect 361690 167 362718 856
rect 362886 167 363914 856
rect 364082 167 365110 856
rect 365278 167 366306 856
rect 366474 167 367502 856
rect 367670 167 368698 856
rect 368866 167 369894 856
rect 370062 167 371090 856
rect 371258 167 372286 856
rect 372454 167 373482 856
rect 373650 167 374678 856
rect 374846 167 375874 856
rect 376042 167 377070 856
rect 377238 167 378266 856
rect 378434 167 379462 856
rect 379630 167 380658 856
rect 380826 167 381854 856
rect 382022 167 383050 856
rect 383218 167 384246 856
rect 384414 167 385442 856
rect 385610 167 386638 856
rect 386806 167 387834 856
rect 388002 167 389030 856
rect 389198 167 390226 856
rect 390394 167 391422 856
rect 391590 167 392618 856
rect 392786 167 393814 856
rect 393982 167 395010 856
rect 395178 167 396206 856
rect 396374 167 397402 856
rect 397570 167 398598 856
rect 398766 167 399794 856
rect 399962 167 400990 856
rect 401158 167 402186 856
rect 402354 167 403382 856
rect 403550 167 404578 856
rect 404746 167 405774 856
rect 405942 167 406970 856
rect 407138 167 408166 856
rect 408334 167 409362 856
rect 409530 167 410558 856
rect 410726 167 411754 856
rect 411922 167 412950 856
rect 413118 167 414146 856
rect 414314 167 415342 856
rect 415510 167 416538 856
rect 416706 167 417734 856
rect 417902 167 418930 856
rect 419098 167 420126 856
rect 420294 167 421322 856
rect 421490 167 422518 856
rect 422686 167 423714 856
rect 423882 167 424910 856
rect 425078 167 426106 856
rect 426274 167 427302 856
rect 427470 167 428498 856
rect 428666 167 429694 856
rect 429862 167 430890 856
rect 431058 167 432086 856
rect 432254 167 433282 856
rect 433450 167 434478 856
rect 434646 167 435674 856
rect 435842 167 436870 856
rect 437038 167 438066 856
rect 438234 167 439262 856
rect 439430 167 440458 856
rect 440626 167 441654 856
rect 441822 167 442850 856
rect 443018 167 444046 856
rect 444214 167 445242 856
rect 445410 167 446438 856
rect 446606 167 447634 856
rect 447802 167 448830 856
rect 448998 167 450026 856
rect 450194 167 451222 856
rect 451390 167 452418 856
rect 452586 167 453614 856
rect 453782 167 454810 856
rect 454978 167 456006 856
rect 456174 167 457202 856
rect 457370 167 458398 856
rect 458566 167 459594 856
rect 459762 167 460790 856
rect 460958 167 461986 856
rect 462154 167 463182 856
rect 463350 167 464378 856
rect 464546 167 465574 856
rect 465742 167 466770 856
rect 466938 167 467966 856
rect 468134 167 469162 856
rect 469330 167 470358 856
rect 470526 167 471554 856
rect 471722 167 472750 856
rect 472918 167 473946 856
rect 474114 167 475142 856
rect 475310 167 476338 856
rect 476506 167 477534 856
rect 477702 167 478730 856
rect 478898 167 479926 856
rect 480094 167 481122 856
rect 481290 167 482318 856
rect 482486 167 483514 856
rect 483682 167 484710 856
rect 484878 167 485906 856
rect 486074 167 487102 856
rect 487270 167 488298 856
rect 488466 167 489494 856
rect 489662 167 490690 856
rect 490858 167 491886 856
rect 492054 167 493082 856
rect 493250 167 494278 856
rect 494446 167 495474 856
rect 495642 167 496670 856
rect 496838 167 497866 856
rect 498034 167 499062 856
rect 499230 167 500258 856
rect 500426 167 501454 856
rect 501622 167 502650 856
rect 502818 167 503846 856
rect 504014 167 505042 856
rect 505210 167 506238 856
rect 506406 167 507434 856
rect 507602 167 508630 856
rect 508798 167 509826 856
rect 509994 167 511022 856
rect 511190 167 512218 856
rect 512386 167 513414 856
rect 513582 167 514610 856
rect 514778 167 515806 856
rect 515974 167 517002 856
rect 517170 167 518198 856
rect 518366 167 519394 856
rect 519562 167 520590 856
rect 520758 167 521786 856
rect 521954 167 522982 856
rect 523150 167 524178 856
rect 524346 167 525374 856
rect 525542 167 526570 856
rect 526738 167 527766 856
rect 527934 167 528962 856
rect 529130 167 530158 856
rect 530326 167 531354 856
rect 531522 167 532550 856
rect 532718 167 533746 856
rect 533914 167 534942 856
rect 535110 167 536138 856
rect 536306 167 537334 856
rect 537502 167 538530 856
rect 538698 167 539726 856
rect 539894 167 540922 856
rect 541090 167 542118 856
rect 542286 167 543314 856
rect 543482 167 544510 856
rect 544678 167 545706 856
rect 545874 167 546902 856
rect 547070 167 548098 856
rect 548266 167 549294 856
rect 549462 167 550490 856
rect 550658 167 551686 856
rect 551854 167 552882 856
rect 553050 167 554078 856
rect 554246 167 555274 856
rect 555442 167 556470 856
rect 556638 167 557666 856
rect 557834 167 558862 856
rect 559030 167 560058 856
rect 560226 167 561254 856
rect 561422 167 562450 856
rect 562618 167 563646 856
rect 563814 167 564842 856
rect 565010 167 566038 856
rect 566206 167 567234 856
rect 567402 167 568430 856
rect 568598 167 569626 856
rect 569794 167 570822 856
rect 570990 167 572018 856
rect 572186 167 573214 856
rect 573382 167 574410 856
rect 574578 167 575606 856
rect 575774 167 576802 856
rect 576970 167 577998 856
rect 578166 167 579194 856
rect 579362 167 580390 856
rect 580558 167 581586 856
rect 581754 167 582782 856
rect 582950 167 583978 856
rect 584146 167 585174 856
rect 585342 167 586370 856
rect 586538 167 587566 856
rect 587734 167 588762 856
rect 588930 167 589958 856
rect 590126 167 591154 856
rect 591322 167 592350 856
rect 592518 167 593546 856
rect 593714 167 594742 856
rect 594910 167 599546 856
<< metal3 >>
rect 600400 709520 601200 709640
rect 0 708024 800 708144
rect 600400 693608 601200 693728
rect 0 691024 800 691144
rect 600400 677696 601200 677816
rect 0 674024 800 674144
rect 600400 661784 601200 661904
rect 0 657024 800 657144
rect 600400 645872 601200 645992
rect 0 640024 800 640144
rect 600400 629960 601200 630080
rect 0 623024 800 623144
rect 600400 614048 601200 614168
rect 0 606024 800 606144
rect 600400 598136 601200 598256
rect 0 589024 800 589144
rect 600400 582224 601200 582344
rect 0 572024 800 572144
rect 600400 566312 601200 566432
rect 0 555024 800 555144
rect 600400 550400 601200 550520
rect 0 538024 800 538144
rect 600400 534488 601200 534608
rect 0 521024 800 521144
rect 600400 518576 601200 518696
rect 0 504024 800 504144
rect 600400 502664 601200 502784
rect 0 487024 800 487144
rect 600400 486752 601200 486872
rect 600400 470840 601200 470960
rect 0 470024 800 470144
rect 600400 454928 601200 455048
rect 0 453024 800 453144
rect 600400 439016 601200 439136
rect 0 436024 800 436144
rect 600400 423104 601200 423224
rect 0 419024 800 419144
rect 600400 407192 601200 407312
rect 0 402024 800 402144
rect 600400 391280 601200 391400
rect 0 385024 800 385144
rect 600400 375368 601200 375488
rect 0 368024 800 368144
rect 600400 359456 601200 359576
rect 0 351024 800 351144
rect 600400 343544 601200 343664
rect 0 334024 800 334144
rect 600400 327632 601200 327752
rect 0 317024 800 317144
rect 600400 311720 601200 311840
rect 0 300024 800 300144
rect 600400 295808 601200 295928
rect 0 283024 800 283144
rect 600400 279896 601200 280016
rect 0 266024 800 266144
rect 600400 263984 601200 264104
rect 0 249024 800 249144
rect 600400 248072 601200 248192
rect 0 232024 800 232144
rect 600400 232160 601200 232280
rect 600400 216248 601200 216368
rect 0 215024 800 215144
rect 600400 200336 601200 200456
rect 0 198024 800 198144
rect 600400 184424 601200 184544
rect 0 181024 800 181144
rect 600400 168512 601200 168632
rect 0 164024 800 164144
rect 600400 152600 601200 152720
rect 0 147024 800 147144
rect 600400 136688 601200 136808
rect 0 130024 800 130144
rect 600400 120776 601200 120896
rect 0 113024 800 113144
rect 600400 104864 601200 104984
rect 0 96024 800 96144
rect 600400 88952 601200 89072
rect 0 79024 800 79144
rect 600400 73040 601200 73160
rect 0 62024 800 62144
rect 600400 57128 601200 57248
rect 0 45024 800 45144
rect 600400 41216 601200 41336
rect 0 28024 800 28144
rect 600400 25304 601200 25424
rect 0 11024 800 11144
rect 600400 9392 601200 9512
<< obsm3 >>
rect 800 709720 600400 717025
rect 800 709440 600320 709720
rect 800 708224 600400 709440
rect 880 707944 600400 708224
rect 800 693808 600400 707944
rect 800 693528 600320 693808
rect 800 691224 600400 693528
rect 880 690944 600400 691224
rect 800 677896 600400 690944
rect 800 677616 600320 677896
rect 800 674224 600400 677616
rect 880 673944 600400 674224
rect 800 661984 600400 673944
rect 800 661704 600320 661984
rect 800 657224 600400 661704
rect 880 656944 600400 657224
rect 800 646072 600400 656944
rect 800 645792 600320 646072
rect 800 640224 600400 645792
rect 880 639944 600400 640224
rect 800 630160 600400 639944
rect 800 629880 600320 630160
rect 800 623224 600400 629880
rect 880 622944 600400 623224
rect 800 614248 600400 622944
rect 800 613968 600320 614248
rect 800 606224 600400 613968
rect 880 605944 600400 606224
rect 800 598336 600400 605944
rect 800 598056 600320 598336
rect 800 589224 600400 598056
rect 880 588944 600400 589224
rect 800 582424 600400 588944
rect 800 582144 600320 582424
rect 800 572224 600400 582144
rect 880 571944 600400 572224
rect 800 566512 600400 571944
rect 800 566232 600320 566512
rect 800 555224 600400 566232
rect 880 554944 600400 555224
rect 800 550600 600400 554944
rect 800 550320 600320 550600
rect 800 538224 600400 550320
rect 880 537944 600400 538224
rect 800 534688 600400 537944
rect 800 534408 600320 534688
rect 800 521224 600400 534408
rect 880 520944 600400 521224
rect 800 518776 600400 520944
rect 800 518496 600320 518776
rect 800 504224 600400 518496
rect 880 503944 600400 504224
rect 800 502864 600400 503944
rect 800 502584 600320 502864
rect 800 487224 600400 502584
rect 880 486952 600400 487224
rect 880 486944 600320 486952
rect 800 486672 600320 486944
rect 800 471040 600400 486672
rect 800 470760 600320 471040
rect 800 470224 600400 470760
rect 880 469944 600400 470224
rect 800 455128 600400 469944
rect 800 454848 600320 455128
rect 800 453224 600400 454848
rect 880 452944 600400 453224
rect 800 439216 600400 452944
rect 800 438936 600320 439216
rect 800 436224 600400 438936
rect 880 435944 600400 436224
rect 800 423304 600400 435944
rect 800 423024 600320 423304
rect 800 419224 600400 423024
rect 880 418944 600400 419224
rect 800 407392 600400 418944
rect 800 407112 600320 407392
rect 800 402224 600400 407112
rect 880 401944 600400 402224
rect 800 391480 600400 401944
rect 800 391200 600320 391480
rect 800 385224 600400 391200
rect 880 384944 600400 385224
rect 800 375568 600400 384944
rect 800 375288 600320 375568
rect 800 368224 600400 375288
rect 880 367944 600400 368224
rect 800 359656 600400 367944
rect 800 359376 600320 359656
rect 800 351224 600400 359376
rect 880 350944 600400 351224
rect 800 343744 600400 350944
rect 800 343464 600320 343744
rect 800 334224 600400 343464
rect 880 333944 600400 334224
rect 800 327832 600400 333944
rect 800 327552 600320 327832
rect 800 317224 600400 327552
rect 880 316944 600400 317224
rect 800 311920 600400 316944
rect 800 311640 600320 311920
rect 800 300224 600400 311640
rect 880 299944 600400 300224
rect 800 296008 600400 299944
rect 800 295728 600320 296008
rect 800 283224 600400 295728
rect 880 282944 600400 283224
rect 800 280096 600400 282944
rect 800 279816 600320 280096
rect 800 266224 600400 279816
rect 880 265944 600400 266224
rect 800 264184 600400 265944
rect 800 263904 600320 264184
rect 800 249224 600400 263904
rect 880 248944 600400 249224
rect 800 248272 600400 248944
rect 800 247992 600320 248272
rect 800 232360 600400 247992
rect 800 232224 600320 232360
rect 880 232080 600320 232224
rect 880 231944 600400 232080
rect 800 216448 600400 231944
rect 800 216168 600320 216448
rect 800 215224 600400 216168
rect 880 214944 600400 215224
rect 800 200536 600400 214944
rect 800 200256 600320 200536
rect 800 198224 600400 200256
rect 880 197944 600400 198224
rect 800 184624 600400 197944
rect 800 184344 600320 184624
rect 800 181224 600400 184344
rect 880 180944 600400 181224
rect 800 168712 600400 180944
rect 800 168432 600320 168712
rect 800 164224 600400 168432
rect 880 163944 600400 164224
rect 800 152800 600400 163944
rect 800 152520 600320 152800
rect 800 147224 600400 152520
rect 880 146944 600400 147224
rect 800 136888 600400 146944
rect 800 136608 600320 136888
rect 800 130224 600400 136608
rect 880 129944 600400 130224
rect 800 120976 600400 129944
rect 800 120696 600320 120976
rect 800 113224 600400 120696
rect 880 112944 600400 113224
rect 800 105064 600400 112944
rect 800 104784 600320 105064
rect 800 96224 600400 104784
rect 880 95944 600400 96224
rect 800 89152 600400 95944
rect 800 88872 600320 89152
rect 800 79224 600400 88872
rect 880 78944 600400 79224
rect 800 73240 600400 78944
rect 800 72960 600320 73240
rect 800 62224 600400 72960
rect 880 61944 600400 62224
rect 800 57328 600400 61944
rect 800 57048 600320 57328
rect 800 45224 600400 57048
rect 880 44944 600400 45224
rect 800 41416 600400 44944
rect 800 41136 600320 41416
rect 800 28224 600400 41136
rect 880 27944 600400 28224
rect 800 25504 600400 27944
rect 800 25224 600320 25504
rect 800 11224 600400 25224
rect 880 10944 600400 11224
rect 800 9592 600400 10944
rect 800 9312 600320 9592
rect 800 171 600400 9312
<< metal4 >>
rect -1076 -4 -756 719172
rect -416 656 -96 718512
rect 2568 -4 6168 719172
rect 7676 580944 11276 706160
rect 17928 705200 21528 719172
rect 33288 705200 36888 719172
rect 48648 705200 52248 719172
rect 64008 705200 67608 719172
rect 79368 705200 82968 719172
rect 94728 705200 98328 719172
rect 110088 705200 113688 719172
rect 125448 705200 129048 719172
rect 140808 705200 144408 719172
rect 156168 705200 159768 719172
rect 171528 705200 175128 719172
rect 186888 705200 190488 719172
rect 7676 440592 11276 565808
rect 17928 565400 21528 581200
rect 33288 565400 36888 581200
rect 48648 565400 52248 581200
rect 64008 565400 67608 581200
rect 79368 565400 82968 581200
rect 94728 565400 98328 581200
rect 110088 565400 113688 581200
rect 125448 565400 129048 581200
rect 140808 565400 144408 581200
rect 156168 565400 159768 581200
rect 171528 565400 175128 581200
rect 186888 565400 190488 581200
rect 7676 301328 11276 426544
rect 17928 425600 21528 441400
rect 33288 425600 36888 441400
rect 48648 425600 52248 441400
rect 64008 425600 67608 441400
rect 79368 425600 82968 441400
rect 94728 425600 98328 441400
rect 110088 425600 113688 441400
rect 125448 425600 129048 441400
rect 140808 425600 144408 441400
rect 156168 425600 159768 441400
rect 171528 425600 175128 441400
rect 186888 425600 190488 441400
rect 7676 160976 11276 286192
rect 17928 285800 21528 301600
rect 33288 285800 36888 301600
rect 48648 285800 52248 301600
rect 64008 285800 67608 301600
rect 79368 285800 82968 301600
rect 94728 285800 98328 301600
rect 110088 285800 113688 301600
rect 125448 285800 129048 301600
rect 140808 285800 144408 301600
rect 156168 285800 159768 301600
rect 171528 285800 175128 301600
rect 186888 285800 190488 301600
rect 7676 19124 11276 146928
rect 17928 146000 21528 161800
rect 33288 146000 36888 161800
rect 48648 146000 52248 161800
rect 64008 146000 67608 161800
rect 79368 146000 82968 161800
rect 94728 146000 98328 161800
rect 110088 146000 113688 161800
rect 125448 146000 129048 161800
rect 140808 146000 144408 161800
rect 156168 146000 159768 161800
rect 171528 146000 175128 161800
rect 186888 146000 190488 161800
rect 17928 -4 21528 22000
rect 33288 -4 36888 22000
rect 48648 -4 52248 22000
rect 64008 -4 67608 22000
rect 79368 -4 82968 22000
rect 94728 -4 98328 22000
rect 110088 -4 113688 22000
rect 125448 -4 129048 22000
rect 140808 -4 144408 22000
rect 156168 -4 159768 22000
rect 171528 -4 175128 22000
rect 186888 -4 190488 22000
rect 202248 -4 205848 719172
rect 206008 580400 207808 705616
rect 217608 705200 221208 719172
rect 232968 705200 236568 719172
rect 248328 705200 251928 719172
rect 263688 705200 267288 719172
rect 279048 705200 282648 719172
rect 294408 705200 298008 719172
rect 309768 705200 313368 719172
rect 325128 705200 328728 719172
rect 340488 705200 344088 719172
rect 355848 705200 359448 719172
rect 371208 705200 374808 719172
rect 386568 705200 390168 719172
rect 206008 441136 207808 569160
rect 217608 565400 221208 581200
rect 232968 565400 236568 581200
rect 248328 565400 251928 581200
rect 263688 565400 267288 581200
rect 279048 565400 282648 581200
rect 294408 565400 298008 581200
rect 309768 565400 313368 581200
rect 325128 565400 328728 581200
rect 340488 565400 344088 581200
rect 355848 565400 359448 581200
rect 371208 565400 374808 581200
rect 386568 565400 390168 581200
rect 394056 580400 395856 706160
rect 396080 580400 397880 706160
rect 401928 705200 405528 719172
rect 417288 705200 420888 719172
rect 432648 705200 436248 719172
rect 448008 705200 451608 719172
rect 463368 705200 466968 719172
rect 478728 705200 482328 719172
rect 494088 705200 497688 719172
rect 509448 705200 513048 719172
rect 524808 705200 528408 719172
rect 540168 705200 543768 719172
rect 555528 705200 559128 719172
rect 570888 705200 574488 719172
rect 206008 300784 207808 426000
rect 217608 425600 221208 441400
rect 232968 425600 236568 441400
rect 248328 425600 251928 441400
rect 263688 425600 267288 441400
rect 279048 425600 282648 441400
rect 294408 425600 298008 441400
rect 309768 425600 313368 441400
rect 325128 425600 328728 441400
rect 340488 425600 344088 441400
rect 355848 425600 359448 441400
rect 371208 425600 374808 441400
rect 386568 425600 390168 441400
rect 394056 440592 395856 569160
rect 396080 440592 397880 566352
rect 401928 565400 405528 581200
rect 417288 565400 420888 581200
rect 432648 565400 436248 581200
rect 448008 565400 451608 581200
rect 463368 565400 466968 581200
rect 478728 565400 482328 581200
rect 494088 565400 497688 581200
rect 509448 565400 513048 581200
rect 524808 565400 528408 581200
rect 540168 565400 543768 581200
rect 555528 565400 559128 581200
rect 570888 565400 574488 581200
rect 206008 161520 207808 286736
rect 217608 285800 221208 301600
rect 232968 285800 236568 301600
rect 248328 285800 251928 301600
rect 263688 285800 267288 301600
rect 279048 285800 282648 301600
rect 294408 285800 298008 301600
rect 309768 285800 313368 301600
rect 325128 285800 328728 301600
rect 340488 285800 344088 301600
rect 355848 285800 359448 301600
rect 371208 285800 374808 301600
rect 386568 285800 390168 301600
rect 394056 300784 395856 426544
rect 396080 300784 397880 426544
rect 401928 425600 405528 441400
rect 417288 425600 420888 441400
rect 432648 425600 436248 441400
rect 448008 425600 451608 441400
rect 463368 425600 466968 441400
rect 478728 425600 482328 441400
rect 494088 425600 497688 441400
rect 509448 425600 513048 441400
rect 524808 425600 528408 441400
rect 540168 425600 543768 441400
rect 555528 425600 559128 441400
rect 570888 425600 574488 441400
rect 206008 21168 207808 146384
rect 217608 146000 221208 161800
rect 232968 146000 236568 161800
rect 248328 146000 251928 161800
rect 263688 146000 267288 161800
rect 279048 146000 282648 161800
rect 294408 146000 298008 161800
rect 309768 146000 313368 161800
rect 325128 146000 328728 161800
rect 340488 146000 344088 161800
rect 355848 146000 359448 161800
rect 371208 146000 374808 161800
rect 386568 146000 390168 161800
rect 394056 160976 395856 286736
rect 396080 160976 397880 286736
rect 401928 285800 405528 301600
rect 417288 285800 420888 301600
rect 432648 285800 436248 301600
rect 448008 285800 451608 301600
rect 463368 285800 466968 301600
rect 478728 285800 482328 301600
rect 494088 285800 497688 301600
rect 509448 285800 513048 301600
rect 524808 285800 528408 301600
rect 540168 285800 543768 301600
rect 555528 285800 559128 301600
rect 570888 285800 574488 301600
rect 217608 -4 221208 22000
rect 232968 -4 236568 22000
rect 248328 -4 251928 22000
rect 263688 -4 267288 22000
rect 279048 -4 282648 22000
rect 294408 -4 298008 22000
rect 309768 -4 313368 22000
rect 325128 -4 328728 22000
rect 340488 -4 344088 22000
rect 355848 -4 359448 22000
rect 371208 -4 374808 22000
rect 386568 -4 390168 22000
rect 394056 21168 395856 146928
rect 396080 19124 397880 146928
rect 401928 146000 405528 161800
rect 417288 146000 420888 161800
rect 432648 146000 436248 161800
rect 448008 146000 451608 161800
rect 463368 146000 466968 161800
rect 478728 146000 482328 161800
rect 494088 146000 497688 161800
rect 509448 146000 513048 161800
rect 524808 146000 528408 161800
rect 540168 146000 543768 161800
rect 555528 146000 559128 161800
rect 570888 146000 574488 161800
rect 401928 -4 405528 22000
rect 417288 -4 420888 22000
rect 432648 -4 436248 22000
rect 448008 -4 451608 22000
rect 463368 -4 466968 22000
rect 478728 -4 482328 22000
rect 494088 -4 497688 22000
rect 509448 -4 513048 22000
rect 524808 -4 528408 22000
rect 540168 -4 543768 22000
rect 555528 -4 559128 22000
rect 570888 -4 574488 22000
rect 586248 -4 589848 719172
rect 594084 580944 597684 706160
rect 594084 440592 597684 565808
rect 594084 301328 597684 426544
rect 594084 160976 597684 286192
rect 594084 19124 597684 146928
rect 601224 656 601544 718512
rect 601884 -4 602204 719172
<< obsm4 >>
rect 2182 579 2488 716685
rect 6248 706240 17848 716685
rect 6248 580864 7596 706240
rect 11356 705120 17848 706240
rect 21608 705120 33208 716685
rect 36968 705120 48568 716685
rect 52328 705120 63928 716685
rect 67688 705120 79288 716685
rect 83048 705120 94648 716685
rect 98408 705120 110008 716685
rect 113768 705120 125368 716685
rect 129128 705120 140728 716685
rect 144488 705120 156088 716685
rect 159848 705120 171448 716685
rect 175208 705120 186808 716685
rect 190568 705120 202168 716685
rect 11356 581280 202168 705120
rect 11356 580864 17848 581280
rect 6248 565888 17848 580864
rect 6248 440512 7596 565888
rect 11356 565320 17848 565888
rect 21608 565320 33208 581280
rect 36968 565320 48568 581280
rect 52328 565320 63928 581280
rect 67688 565320 79288 581280
rect 83048 565320 94648 581280
rect 98408 565320 110008 581280
rect 113768 565320 125368 581280
rect 129128 565320 140728 581280
rect 144488 565320 156088 581280
rect 159848 565320 171448 581280
rect 175208 565320 186808 581280
rect 190568 565320 202168 581280
rect 11356 441480 202168 565320
rect 11356 440512 17848 441480
rect 6248 426624 17848 440512
rect 6248 301248 7596 426624
rect 11356 425520 17848 426624
rect 21608 425520 33208 441480
rect 36968 425520 48568 441480
rect 52328 425520 63928 441480
rect 67688 425520 79288 441480
rect 83048 425520 94648 441480
rect 98408 425520 110008 441480
rect 113768 425520 125368 441480
rect 129128 425520 140728 441480
rect 144488 425520 156088 441480
rect 159848 425520 171448 441480
rect 175208 425520 186808 441480
rect 190568 425520 202168 441480
rect 11356 301680 202168 425520
rect 11356 301248 17848 301680
rect 6248 286272 17848 301248
rect 6248 160896 7596 286272
rect 11356 285720 17848 286272
rect 21608 285720 33208 301680
rect 36968 285720 48568 301680
rect 52328 285720 63928 301680
rect 67688 285720 79288 301680
rect 83048 285720 94648 301680
rect 98408 285720 110008 301680
rect 113768 285720 125368 301680
rect 129128 285720 140728 301680
rect 144488 285720 156088 301680
rect 159848 285720 171448 301680
rect 175208 285720 186808 301680
rect 190568 285720 202168 301680
rect 11356 161880 202168 285720
rect 11356 160896 17848 161880
rect 6248 147008 17848 160896
rect 6248 19044 7596 147008
rect 11356 145920 17848 147008
rect 21608 145920 33208 161880
rect 36968 145920 48568 161880
rect 52328 145920 63928 161880
rect 67688 145920 79288 161880
rect 83048 145920 94648 161880
rect 98408 145920 110008 161880
rect 113768 145920 125368 161880
rect 129128 145920 140728 161880
rect 144488 145920 156088 161880
rect 159848 145920 171448 161880
rect 175208 145920 186808 161880
rect 190568 145920 202168 161880
rect 11356 22080 202168 145920
rect 11356 19044 17848 22080
rect 6248 579 17848 19044
rect 21608 579 33208 22080
rect 36968 579 48568 22080
rect 52328 579 63928 22080
rect 67688 579 79288 22080
rect 83048 579 94648 22080
rect 98408 579 110008 22080
rect 113768 579 125368 22080
rect 129128 579 140728 22080
rect 144488 579 156088 22080
rect 159848 579 171448 22080
rect 175208 579 186808 22080
rect 190568 579 202168 22080
rect 205928 705696 217528 716685
rect 207888 705120 217528 705696
rect 221288 705120 232888 716685
rect 236648 705120 248248 716685
rect 252008 705120 263608 716685
rect 267368 705120 278968 716685
rect 282728 705120 294328 716685
rect 298088 705120 309688 716685
rect 313448 705120 325048 716685
rect 328808 705120 340408 716685
rect 344168 705120 355768 716685
rect 359528 705120 371128 716685
rect 374888 705120 386488 716685
rect 390248 706240 401848 716685
rect 390248 705120 393976 706240
rect 207888 581280 393976 705120
rect 207888 580320 217528 581280
rect 205928 569240 217528 580320
rect 207888 565320 217528 569240
rect 221288 565320 232888 581280
rect 236648 565320 248248 581280
rect 252008 565320 263608 581280
rect 267368 565320 278968 581280
rect 282728 565320 294328 581280
rect 298088 565320 309688 581280
rect 313448 565320 325048 581280
rect 328808 565320 340408 581280
rect 344168 565320 355768 581280
rect 359528 565320 371128 581280
rect 374888 565320 386488 581280
rect 390248 580320 393976 581280
rect 395936 580320 396000 706240
rect 397960 705120 401848 706240
rect 405608 705120 417208 716685
rect 420968 705120 432568 716685
rect 436328 705120 447928 716685
rect 451688 705120 463288 716685
rect 467048 705120 478648 716685
rect 482408 705120 494008 716685
rect 497768 705120 509368 716685
rect 513128 705120 524728 716685
rect 528488 705120 540088 716685
rect 543848 705120 555448 716685
rect 559208 705120 570808 716685
rect 574568 705120 586168 716685
rect 397960 581280 586168 705120
rect 397960 580320 401848 581280
rect 390248 569240 401848 580320
rect 390248 565320 393976 569240
rect 207888 441480 393976 565320
rect 207888 441056 217528 441480
rect 205928 426080 217528 441056
rect 207888 425520 217528 426080
rect 221288 425520 232888 441480
rect 236648 425520 248248 441480
rect 252008 425520 263608 441480
rect 267368 425520 278968 441480
rect 282728 425520 294328 441480
rect 298088 425520 309688 441480
rect 313448 425520 325048 441480
rect 328808 425520 340408 441480
rect 344168 425520 355768 441480
rect 359528 425520 371128 441480
rect 374888 425520 386488 441480
rect 390248 440512 393976 441480
rect 395936 566432 401848 569240
rect 395936 440512 396000 566432
rect 397960 565320 401848 566432
rect 405608 565320 417208 581280
rect 420968 565320 432568 581280
rect 436328 565320 447928 581280
rect 451688 565320 463288 581280
rect 467048 565320 478648 581280
rect 482408 565320 494008 581280
rect 497768 565320 509368 581280
rect 513128 565320 524728 581280
rect 528488 565320 540088 581280
rect 543848 565320 555448 581280
rect 559208 565320 570808 581280
rect 574568 565320 586168 581280
rect 397960 441480 586168 565320
rect 397960 440512 401848 441480
rect 390248 426624 401848 440512
rect 390248 425520 393976 426624
rect 207888 301680 393976 425520
rect 207888 300704 217528 301680
rect 205928 286816 217528 300704
rect 207888 285720 217528 286816
rect 221288 285720 232888 301680
rect 236648 285720 248248 301680
rect 252008 285720 263608 301680
rect 267368 285720 278968 301680
rect 282728 285720 294328 301680
rect 298088 285720 309688 301680
rect 313448 285720 325048 301680
rect 328808 285720 340408 301680
rect 344168 285720 355768 301680
rect 359528 285720 371128 301680
rect 374888 285720 386488 301680
rect 390248 300704 393976 301680
rect 395936 300704 396000 426624
rect 397960 425520 401848 426624
rect 405608 425520 417208 441480
rect 420968 425520 432568 441480
rect 436328 425520 447928 441480
rect 451688 425520 463288 441480
rect 467048 425520 478648 441480
rect 482408 425520 494008 441480
rect 497768 425520 509368 441480
rect 513128 425520 524728 441480
rect 528488 425520 540088 441480
rect 543848 425520 555448 441480
rect 559208 425520 570808 441480
rect 574568 425520 586168 441480
rect 397960 301680 586168 425520
rect 397960 300704 401848 301680
rect 390248 286816 401848 300704
rect 390248 285720 393976 286816
rect 207888 161880 393976 285720
rect 207888 161440 217528 161880
rect 205928 146464 217528 161440
rect 207888 145920 217528 146464
rect 221288 145920 232888 161880
rect 236648 145920 248248 161880
rect 252008 145920 263608 161880
rect 267368 145920 278968 161880
rect 282728 145920 294328 161880
rect 298088 145920 309688 161880
rect 313448 145920 325048 161880
rect 328808 145920 340408 161880
rect 344168 145920 355768 161880
rect 359528 145920 371128 161880
rect 374888 145920 386488 161880
rect 390248 160896 393976 161880
rect 395936 160896 396000 286816
rect 397960 285720 401848 286816
rect 405608 285720 417208 301680
rect 420968 285720 432568 301680
rect 436328 285720 447928 301680
rect 451688 285720 463288 301680
rect 467048 285720 478648 301680
rect 482408 285720 494008 301680
rect 497768 285720 509368 301680
rect 513128 285720 524728 301680
rect 528488 285720 540088 301680
rect 543848 285720 555448 301680
rect 559208 285720 570808 301680
rect 574568 285720 586168 301680
rect 397960 161880 586168 285720
rect 397960 160896 401848 161880
rect 390248 147008 401848 160896
rect 390248 145920 393976 147008
rect 207888 22080 393976 145920
rect 207888 21088 217528 22080
rect 205928 579 217528 21088
rect 221288 579 232888 22080
rect 236648 579 248248 22080
rect 252008 579 263608 22080
rect 267368 579 278968 22080
rect 282728 579 294328 22080
rect 298088 579 309688 22080
rect 313448 579 325048 22080
rect 328808 579 340408 22080
rect 344168 579 355768 22080
rect 359528 579 371128 22080
rect 374888 579 386488 22080
rect 390248 21088 393976 22080
rect 395936 21088 396000 147008
rect 390248 19044 396000 21088
rect 397960 145920 401848 147008
rect 405608 145920 417208 161880
rect 420968 145920 432568 161880
rect 436328 145920 447928 161880
rect 451688 145920 463288 161880
rect 467048 145920 478648 161880
rect 482408 145920 494008 161880
rect 497768 145920 509368 161880
rect 513128 145920 524728 161880
rect 528488 145920 540088 161880
rect 543848 145920 555448 161880
rect 559208 145920 570808 161880
rect 574568 145920 586168 161880
rect 397960 22080 586168 145920
rect 397960 19044 401848 22080
rect 390248 579 401848 19044
rect 405608 579 417208 22080
rect 420968 579 432568 22080
rect 436328 579 447928 22080
rect 451688 579 463288 22080
rect 467048 579 478648 22080
rect 482408 579 494008 22080
rect 497768 579 509368 22080
rect 513128 579 524728 22080
rect 528488 579 540088 22080
rect 543848 579 555448 22080
rect 559208 579 570808 22080
rect 574568 579 586168 22080
rect 589928 706240 598026 716685
rect 589928 580864 594004 706240
rect 597764 580864 598026 706240
rect 589928 565888 598026 580864
rect 589928 440512 594004 565888
rect 597764 440512 598026 565888
rect 589928 426624 598026 440512
rect 589928 301248 594004 426624
rect 597764 301248 598026 426624
rect 589928 286272 598026 301248
rect 589928 160896 594004 286272
rect 597764 160896 598026 286272
rect 589928 147008 598026 160896
rect 589928 19044 594004 147008
rect 597764 19044 598026 147008
rect 589928 579 598026 19044
<< metal5 >>
rect -1076 718852 602204 719172
rect -416 718192 601544 718512
rect -1076 708434 602204 711834
rect -1076 693116 602204 696516
rect -1076 677798 602204 681198
rect -1076 662480 602204 665880
rect -1076 647162 602204 650562
rect -1076 631844 602204 635244
rect -1076 616526 602204 619926
rect -1076 601208 602204 604608
rect -1076 585890 602204 589290
rect -1076 570572 602204 573972
rect 2568 565760 589848 569160
rect -1076 555254 602204 558654
rect -1076 539936 602204 543336
rect -1076 524618 602204 528018
rect -1076 509300 602204 512700
rect -1076 493982 602204 497382
rect -1076 478664 602204 482064
rect -1076 463346 602204 466746
rect -1076 448028 602204 451428
rect -1076 432710 602204 436110
rect 1056 427720 600072 431120
rect -1076 417392 602204 420792
rect -1076 402074 602204 405474
rect -1076 386756 602204 390156
rect -1076 371438 602204 374838
rect -1076 356120 602204 359520
rect -1076 340802 602204 344202
rect -1076 325484 602204 328884
rect -1076 310166 602204 313566
rect -1076 294848 602204 298248
rect 2568 288320 589848 291720
rect -1076 279530 602204 282930
rect -1076 264212 602204 267612
rect -1076 248894 602204 252294
rect -1076 233576 602204 236976
rect -1076 218258 602204 221658
rect -1076 202940 602204 206340
rect -1076 187622 602204 191022
rect -1076 172304 602204 175704
rect -1076 156986 602204 160386
rect 1056 152320 600072 155720
rect -1076 141668 602204 145068
rect -1076 126350 602204 129750
rect -1076 111032 602204 114432
rect -1076 95714 602204 99114
rect -1076 80396 602204 83796
rect -1076 65078 602204 68478
rect -1076 49760 602204 53160
rect -1076 34442 602204 37842
rect -1076 19124 602204 22524
rect -1076 3806 602204 7206
rect -416 656 601544 976
rect -1076 -4 602204 316
<< obsm5 >>
rect 2140 650882 598068 655340
rect 2140 635564 598068 646842
rect 2140 620246 598068 631524
rect 2140 604928 598068 616206
rect 2140 589610 598068 600888
rect 2140 574292 598068 585570
rect 2140 569480 598068 570252
rect 2140 565440 2248 569480
rect 590168 565440 598068 569480
rect 2140 558974 598068 565440
rect 2140 543656 598068 554934
rect 2140 528338 598068 539616
rect 2140 513020 598068 524298
rect 2140 497702 598068 508980
rect 2140 482384 598068 493662
rect 2140 467066 598068 478344
rect 2140 451748 598068 463026
rect 2140 436430 598068 447708
rect 2140 431440 598068 432390
rect 2140 421112 598068 427400
rect 2140 405794 598068 417072
rect 2140 390476 598068 401754
rect 2140 375158 598068 386436
rect 2140 359840 598068 371118
rect 2140 344522 598068 355800
rect 2140 329204 598068 340482
rect 2140 313886 598068 325164
rect 2140 298568 598068 309846
rect 2140 292040 598068 294528
rect 2140 288000 2248 292040
rect 590168 288000 598068 292040
rect 2140 283250 598068 288000
rect 2140 267932 598068 279210
rect 2140 252614 598068 263892
rect 2140 237296 598068 248574
rect 2140 221978 598068 233256
rect 2140 206660 598068 217938
rect 2140 191342 598068 202620
rect 2140 176024 598068 187302
rect 2140 160706 598068 171984
rect 2140 156040 598068 156666
rect 2140 145388 598068 152000
rect 2140 130070 598068 141348
rect 2140 114752 598068 126030
rect 2140 99434 598068 110712
rect 2140 84116 598068 95394
rect 2140 68798 598068 80076
rect 2140 53480 598068 64758
rect 2140 38162 598068 49440
rect 2140 22844 598068 34122
rect 2140 7526 598068 18804
rect 2140 1540 598068 3486
<< labels >>
rlabel metal3 s 600400 9392 601200 9512 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 600400 486752 601200 486872 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 600400 534488 601200 534608 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 600400 582224 601200 582344 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 600400 629960 601200 630080 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 600400 677696 601200 677816 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 590014 718400 590070 719200 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 523222 718400 523278 719200 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 456430 718400 456486 719200 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 389638 718400 389694 719200 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 322846 718400 322902 719200 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 600400 57128 601200 57248 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 256054 718400 256110 719200 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 189262 718400 189318 719200 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 122470 718400 122526 719200 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 55678 718400 55734 719200 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 708024 800 708144 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 657024 800 657144 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 606024 800 606144 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 555024 800 555144 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 504024 800 504144 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 453024 800 453144 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 600400 104864 601200 104984 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 402024 800 402144 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 351024 800 351144 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 300024 800 300144 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 249024 800 249144 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 198024 800 198144 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 147024 800 147144 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 600400 152600 601200 152720 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 600400 200336 601200 200456 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 600400 248072 601200 248192 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 600400 295808 601200 295928 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 600400 343544 601200 343664 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 600400 391280 601200 391400 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 600400 439016 601200 439136 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 600400 41216 601200 41336 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 600400 518576 601200 518696 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 600400 566312 601200 566432 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 600400 614048 601200 614168 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 600400 661784 601200 661904 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 600400 709520 601200 709640 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 545486 718400 545542 719200 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 478694 718400 478750 719200 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 411902 718400 411958 719200 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 345110 718400 345166 719200 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 278318 718400 278374 719200 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 600400 88952 601200 89072 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 211526 718400 211582 719200 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 144734 718400 144790 719200 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 77942 718400 77998 719200 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 11150 718400 11206 719200 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 674024 800 674144 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 623024 800 623144 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 572024 800 572144 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 521024 800 521144 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 470024 800 470144 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 419024 800 419144 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 600400 136688 601200 136808 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 368024 800 368144 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 317024 800 317144 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 266024 800 266144 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 215024 800 215144 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 164024 800 164144 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 113024 800 113144 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 11024 800 11144 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 600400 184424 601200 184544 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 600400 232160 601200 232280 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 600400 279896 601200 280016 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 600400 327632 601200 327752 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 600400 375368 601200 375488 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 600400 423104 601200 423224 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 600400 470840 601200 470960 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 600400 25304 601200 25424 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 600400 502664 601200 502784 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 600400 550400 601200 550520 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 600400 598136 601200 598256 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 600400 645872 601200 645992 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 600400 693608 601200 693728 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 567750 718400 567806 719200 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 500958 718400 501014 719200 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 434166 718400 434222 719200 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 367374 718400 367430 719200 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 300582 718400 300638 719200 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 600400 73040 601200 73160 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 233790 718400 233846 719200 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 166998 718400 167054 719200 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 100206 718400 100262 719200 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 33414 718400 33470 719200 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 691024 800 691144 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 640024 800 640144 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 589024 800 589144 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 538024 800 538144 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 487024 800 487144 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 436024 800 436144 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 600400 120776 601200 120896 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 385024 800 385144 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 334024 800 334144 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 283024 800 283144 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 232024 800 232144 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 181024 800 181144 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 130024 800 130144 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 79024 800 79144 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 600400 168512 601200 168632 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 600400 216248 601200 216368 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 600400 263984 601200 264104 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 600400 311720 601200 311840 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 600400 359456 601200 359576 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 600400 407192 601200 407312 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 600400 454928 601200 455048 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 592406 0 592462 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 593602 0 593658 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 594798 0 594854 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 491942 0 491998 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 495530 0 495586 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 499118 0 499174 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 502706 0 502762 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 506294 0 506350 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 509882 0 509938 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 513470 0 513526 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 517058 0 517114 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 520646 0 520702 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 524234 0 524290 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 527822 0 527878 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 531410 0 531466 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 534998 0 535054 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 538586 0 538642 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 542174 0 542230 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 545762 0 545818 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 549350 0 549406 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 552938 0 552994 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 556526 0 556582 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 560114 0 560170 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 563702 0 563758 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 567290 0 567346 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 570878 0 570934 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 574466 0 574522 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 578054 0 578110 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 581642 0 581698 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 585230 0 585286 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 588818 0 588874 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 183374 0 183430 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 190550 0 190606 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 194138 0 194194 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 201314 0 201370 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 204902 0 204958 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 208490 0 208546 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 212078 0 212134 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 215666 0 215722 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 219254 0 219310 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 222842 0 222898 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 226430 0 226486 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 230018 0 230074 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 233606 0 233662 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 237194 0 237250 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 240782 0 240838 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 244370 0 244426 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 247958 0 248014 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 251546 0 251602 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 255134 0 255190 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 258722 0 258778 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 262310 0 262366 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 265898 0 265954 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 269486 0 269542 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 273074 0 273130 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 276662 0 276718 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 280250 0 280306 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 283838 0 283894 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 287426 0 287482 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 291014 0 291070 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 294602 0 294658 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 298190 0 298246 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 301778 0 301834 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 305366 0 305422 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 308954 0 309010 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 312542 0 312598 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 316130 0 316186 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 319718 0 319774 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 323306 0 323362 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 326894 0 326950 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 330482 0 330538 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 334070 0 334126 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 337658 0 337714 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 341246 0 341302 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 344834 0 344890 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 348422 0 348478 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 352010 0 352066 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 355598 0 355654 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 359186 0 359242 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 362774 0 362830 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 366362 0 366418 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 369950 0 370006 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 373538 0 373594 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 377126 0 377182 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 380714 0 380770 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 384302 0 384358 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 387890 0 387946 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 391478 0 391534 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 395066 0 395122 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 398654 0 398710 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 402242 0 402298 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 405830 0 405886 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 409418 0 409474 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 413006 0 413062 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 416594 0 416650 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 420182 0 420238 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 423770 0 423826 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 427358 0 427414 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 430946 0 431002 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 434534 0 434590 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 438122 0 438178 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 441710 0 441766 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 445298 0 445354 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 448886 0 448942 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 452474 0 452530 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 456062 0 456118 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 459650 0 459706 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 463238 0 463294 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 466826 0 466882 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 470414 0 470470 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 474002 0 474058 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 477590 0 477646 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 481178 0 481234 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 484766 0 484822 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 488354 0 488410 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 493138 0 493194 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 496726 0 496782 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 500314 0 500370 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 503902 0 503958 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 507490 0 507546 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 511078 0 511134 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 514666 0 514722 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 518254 0 518310 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 521842 0 521898 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 525430 0 525486 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 170218 0 170274 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 529018 0 529074 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 532606 0 532662 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 536194 0 536250 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 539782 0 539838 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 543370 0 543426 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 546958 0 547014 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 550546 0 550602 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 554134 0 554190 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 557722 0 557778 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 561310 0 561366 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 173806 0 173862 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 564898 0 564954 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 568486 0 568542 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 572074 0 572130 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 575662 0 575718 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 579250 0 579306 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 582838 0 582894 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 586426 0 586482 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 590014 0 590070 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 177394 0 177450 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 180982 0 181038 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 184570 0 184626 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 188158 0 188214 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 191746 0 191802 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 195334 0 195390 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 198922 0 198978 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 202510 0 202566 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 137926 0 137982 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 206098 0 206154 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 209686 0 209742 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 213274 0 213330 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 216862 0 216918 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 220450 0 220506 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 224038 0 224094 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 227626 0 227682 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 231214 0 231270 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 234802 0 234858 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 238390 0 238446 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 141514 0 141570 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 241978 0 242034 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 245566 0 245622 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 249154 0 249210 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 252742 0 252798 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 256330 0 256386 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 259918 0 259974 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 263506 0 263562 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 267094 0 267150 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 270682 0 270738 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 274270 0 274326 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 145102 0 145158 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 277858 0 277914 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 281446 0 281502 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 285034 0 285090 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 288622 0 288678 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 292210 0 292266 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 295798 0 295854 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 299386 0 299442 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 302974 0 303030 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 306562 0 306618 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 310150 0 310206 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 148690 0 148746 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 313738 0 313794 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 317326 0 317382 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 320914 0 320970 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 324502 0 324558 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 328090 0 328146 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 331678 0 331734 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 335266 0 335322 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 338854 0 338910 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 342442 0 342498 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 346030 0 346086 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 349618 0 349674 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 353206 0 353262 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 356794 0 356850 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 360382 0 360438 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 363970 0 364026 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 367558 0 367614 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 371146 0 371202 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 374734 0 374790 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 378322 0 378378 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 381910 0 381966 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 385498 0 385554 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 389086 0 389142 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 392674 0 392730 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 396262 0 396318 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 399850 0 399906 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 403438 0 403494 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 407026 0 407082 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 410614 0 410670 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 414202 0 414258 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 417790 0 417846 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 159454 0 159510 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 421378 0 421434 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 424966 0 425022 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 428554 0 428610 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 432142 0 432198 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 435730 0 435786 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 439318 0 439374 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 442906 0 442962 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 446494 0 446550 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 450082 0 450138 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 453670 0 453726 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 163042 0 163098 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 457258 0 457314 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 460846 0 460902 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 464434 0 464490 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 468022 0 468078 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 471610 0 471666 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 475198 0 475254 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 478786 0 478842 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 482374 0 482430 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 485962 0 486018 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 489550 0 489606 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 166630 0 166686 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 494334 0 494390 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 497922 0 497978 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 501510 0 501566 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 505098 0 505154 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 508686 0 508742 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 512274 0 512330 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 515862 0 515918 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 519450 0 519506 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 523038 0 523094 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 526626 0 526682 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 171414 0 171470 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 530214 0 530270 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 533802 0 533858 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 537390 0 537446 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 540978 0 541034 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 544566 0 544622 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 548154 0 548210 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 551742 0 551798 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 555330 0 555386 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 558918 0 558974 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 562506 0 562562 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 566094 0 566150 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 569682 0 569738 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 573270 0 573326 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 576858 0 576914 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 580446 0 580502 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 584034 0 584090 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 587622 0 587678 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 591210 0 591266 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 178590 0 178646 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 182178 0 182234 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 185766 0 185822 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 189354 0 189410 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 192942 0 192998 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 200118 0 200174 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 203706 0 203762 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 207294 0 207350 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 210882 0 210938 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 214470 0 214526 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 218058 0 218114 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 221646 0 221702 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 225234 0 225290 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 228822 0 228878 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 232410 0 232466 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 235998 0 236054 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 239586 0 239642 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 243174 0 243230 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 246762 0 246818 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 250350 0 250406 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 253938 0 253994 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 257526 0 257582 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 261114 0 261170 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 264702 0 264758 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 268290 0 268346 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 271878 0 271934 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 275466 0 275522 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 279054 0 279110 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 282642 0 282698 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 286230 0 286286 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 289818 0 289874 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 293406 0 293462 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 296994 0 297050 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 300582 0 300638 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 304170 0 304226 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 307758 0 307814 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 311346 0 311402 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 314934 0 314990 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 318522 0 318578 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 322110 0 322166 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 325698 0 325754 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 329286 0 329342 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 332874 0 332930 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 336462 0 336518 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 340050 0 340106 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 343638 0 343694 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 347226 0 347282 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 350814 0 350870 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 354402 0 354458 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 357990 0 358046 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 361578 0 361634 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 365166 0 365222 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 368754 0 368810 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 372342 0 372398 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 375930 0 375986 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 379518 0 379574 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 383106 0 383162 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 386694 0 386750 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 390282 0 390338 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 393870 0 393926 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 397458 0 397514 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 401046 0 401102 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 404634 0 404690 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 408222 0 408278 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 411810 0 411866 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 415398 0 415454 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 418986 0 419042 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 422574 0 422630 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 426162 0 426218 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 429750 0 429806 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 433338 0 433394 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 436926 0 436982 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 440514 0 440570 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 444102 0 444158 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 447690 0 447746 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 451278 0 451334 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 454866 0 454922 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 458454 0 458510 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 462042 0 462098 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 465630 0 465686 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 469218 0 469274 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 472806 0 472862 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 476394 0 476450 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 479982 0 480038 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 483570 0 483626 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 487158 0 487214 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 490746 0 490802 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 167826 0 167882 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s -416 656 -96 718512 4 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -416 656 601544 976 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -416 718192 601544 718512 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 601224 656 601544 718512 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 2568 -4 6168 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 33288 -4 36888 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 33288 146000 36888 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 33288 285800 36888 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 33288 425600 36888 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 33288 565400 36888 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 33288 705200 36888 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 64008 -4 67608 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 64008 146000 67608 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 64008 285800 67608 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 64008 425600 67608 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 64008 565400 67608 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 64008 705200 67608 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 94728 -4 98328 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 94728 146000 98328 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 94728 285800 98328 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 94728 425600 98328 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 94728 565400 98328 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 94728 705200 98328 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 125448 -4 129048 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 125448 146000 129048 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 125448 285800 129048 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 125448 425600 129048 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 125448 565400 129048 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 125448 705200 129048 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 156168 -4 159768 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 156168 146000 159768 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 156168 285800 159768 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 156168 425600 159768 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 156168 565400 159768 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 156168 705200 159768 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 186888 -4 190488 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 186888 146000 190488 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 186888 285800 190488 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 186888 425600 190488 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 186888 565400 190488 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 186888 705200 190488 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 217608 -4 221208 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 217608 146000 221208 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 217608 285800 221208 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 217608 425600 221208 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 217608 565400 221208 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 217608 705200 221208 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 248328 -4 251928 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 248328 146000 251928 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 248328 285800 251928 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 248328 425600 251928 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 248328 565400 251928 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 248328 705200 251928 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 279048 -4 282648 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 279048 146000 282648 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 279048 285800 282648 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 279048 425600 282648 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 279048 565400 282648 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 279048 705200 282648 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 309768 -4 313368 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 309768 146000 313368 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 309768 285800 313368 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 309768 425600 313368 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 309768 565400 313368 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 309768 705200 313368 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 340488 -4 344088 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 340488 146000 344088 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 340488 285800 344088 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 340488 425600 344088 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 340488 565400 344088 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 340488 705200 344088 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 371208 -4 374808 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 371208 146000 374808 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 371208 285800 374808 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 371208 425600 374808 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 371208 565400 374808 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 371208 705200 374808 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 401928 -4 405528 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 401928 146000 405528 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 401928 285800 405528 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 401928 425600 405528 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 401928 565400 405528 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 401928 705200 405528 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 432648 -4 436248 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 432648 146000 436248 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 432648 285800 436248 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 432648 425600 436248 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 432648 565400 436248 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 432648 705200 436248 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 463368 -4 466968 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 463368 146000 466968 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 463368 285800 466968 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 463368 425600 466968 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 463368 565400 466968 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 463368 705200 466968 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 494088 -4 497688 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 494088 146000 497688 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 494088 285800 497688 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 494088 425600 497688 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 494088 565400 497688 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 494088 705200 497688 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 524808 -4 528408 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 524808 146000 528408 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 524808 285800 528408 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 524808 425600 528408 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 524808 565400 528408 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 524808 705200 528408 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 555528 -4 559128 22000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 555528 146000 559128 161800 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 555528 285800 559128 301600 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 555528 425600 559128 441400 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 555528 565400 559128 581200 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 555528 705200 559128 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 586248 -4 589848 719172 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 3806 602204 7206 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 34442 602204 37842 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 65078 602204 68478 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 95714 602204 99114 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 126350 602204 129750 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 156986 602204 160386 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 187622 602204 191022 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 218258 602204 221658 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 248894 602204 252294 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 279530 602204 282930 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 310166 602204 313566 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 340802 602204 344202 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 371438 602204 374838 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 402074 602204 405474 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 432710 602204 436110 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 463346 602204 466746 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 493982 602204 497382 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 524618 602204 528018 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 555254 602204 558654 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 585890 602204 589290 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 616526 602204 619926 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 647162 602204 650562 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 677798 602204 681198 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 708434 602204 711834 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 206008 161520 207808 286736 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 394056 300784 395856 426544 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 206008 21168 207808 146384 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 394056 440592 395856 569160 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 206008 441136 207808 569160 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 394056 21168 395856 146928 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 206008 300784 207808 426000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 394056 160976 395856 286736 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 206008 580400 207808 705616 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 394056 580400 395856 706160 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s 2568 288320 589848 291720 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s 2568 565760 589848 569160 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s -1076 -4 -756 719172 4 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 -4 602204 316 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 718852 602204 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 601884 -4 602204 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 17928 -4 21528 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 17928 146000 21528 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 17928 285800 21528 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 17928 425600 21528 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 17928 565400 21528 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 17928 705200 21528 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 48648 -4 52248 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 48648 146000 52248 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 48648 285800 52248 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 48648 425600 52248 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 48648 565400 52248 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 48648 705200 52248 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 79368 -4 82968 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 79368 146000 82968 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 79368 285800 82968 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 79368 425600 82968 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 79368 565400 82968 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 79368 705200 82968 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 110088 -4 113688 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 110088 146000 113688 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 110088 285800 113688 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 110088 425600 113688 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 110088 565400 113688 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 110088 705200 113688 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 140808 -4 144408 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 140808 146000 144408 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 140808 285800 144408 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 140808 425600 144408 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 140808 565400 144408 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 140808 705200 144408 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 171528 -4 175128 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 171528 146000 175128 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 171528 285800 175128 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 171528 425600 175128 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 171528 565400 175128 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 171528 705200 175128 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 202248 -4 205848 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 232968 -4 236568 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 232968 146000 236568 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 232968 285800 236568 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 232968 425600 236568 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 232968 565400 236568 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 232968 705200 236568 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 263688 -4 267288 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 263688 146000 267288 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 263688 285800 267288 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 263688 425600 267288 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 263688 565400 267288 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 263688 705200 267288 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 294408 -4 298008 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 294408 146000 298008 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 294408 285800 298008 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 294408 425600 298008 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 294408 565400 298008 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 294408 705200 298008 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 325128 -4 328728 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 325128 146000 328728 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 325128 285800 328728 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 325128 425600 328728 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 325128 565400 328728 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 325128 705200 328728 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 355848 -4 359448 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 355848 146000 359448 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 355848 285800 359448 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 355848 425600 359448 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 355848 565400 359448 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 355848 705200 359448 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 386568 -4 390168 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 386568 146000 390168 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 386568 285800 390168 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 386568 425600 390168 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 386568 565400 390168 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 386568 705200 390168 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 417288 -4 420888 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 417288 146000 420888 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 417288 285800 420888 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 417288 425600 420888 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 417288 565400 420888 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 417288 705200 420888 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 448008 -4 451608 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 448008 146000 451608 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 448008 285800 451608 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 448008 425600 451608 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 448008 565400 451608 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 448008 705200 451608 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 478728 -4 482328 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 478728 146000 482328 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 478728 285800 482328 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 478728 425600 482328 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 478728 565400 482328 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 478728 705200 482328 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 509448 -4 513048 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 509448 146000 513048 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 509448 285800 513048 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 509448 425600 513048 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 509448 565400 513048 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 509448 705200 513048 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 540168 -4 543768 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 540168 146000 543768 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 540168 285800 543768 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 540168 425600 543768 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 540168 565400 543768 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 540168 705200 543768 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 570888 -4 574488 22000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 570888 146000 574488 161800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 570888 285800 574488 301600 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 570888 425600 574488 441400 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 570888 565400 574488 581200 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 570888 705200 574488 719172 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 19124 602204 22524 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 49760 602204 53160 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 80396 602204 83796 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 111032 602204 114432 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 141668 602204 145068 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 172304 602204 175704 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 202940 602204 206340 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 233576 602204 236976 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 264212 602204 267612 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 294848 602204 298248 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 325484 602204 328884 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 356120 602204 359520 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 386756 602204 390156 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 417392 602204 420792 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 448028 602204 451428 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 478664 602204 482064 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 509300 602204 512700 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 539936 602204 543336 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 570572 602204 573972 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 601208 602204 604608 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 631844 602204 635244 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 662480 602204 665880 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 693116 602204 696516 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 7676 19124 11276 146928 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 396080 300784 397880 426544 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 594084 440592 597684 565808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 7676 160976 11276 286192 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 396080 440592 397880 566352 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 594084 301328 597684 426544 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 7676 301328 11276 426544 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 396080 19124 397880 146928 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 594084 160976 597684 286192 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 7676 440592 11276 565808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 396080 160976 397880 286736 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 594084 19124 597684 146928 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 7676 580944 11276 706160 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 396080 580400 397880 706160 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 594084 580944 597684 706160 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s 1056 152320 600072 155720 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s 1056 427720 600072 431120 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 6366 0 6422 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 67362 0 67418 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 103242 0 103298 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 110418 0 110474 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 117594 0 117650 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 124770 0 124826 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 128358 0 128414 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 131946 0 132002 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 601200 719200
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 161221008
string GDS_FILE /home/alex/chaos_automaton_Summer_2022/openlane/chaos_automaton/runs/22_08_10_20_05/results/signoff/chaos_automaton.magic.gds
string GDS_START 54138782
<< end >>

