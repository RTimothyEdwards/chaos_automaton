magic
tech sky130B
magscale 1 2
timestamp 1659633024
<< obsli1 >>
rect 1104 2159 178848 177361
<< obsm1 >>
rect 1104 1912 178848 177540
<< metal2 >>
rect 5170 179200 5226 180000
rect 14094 179200 14150 180000
rect 23018 179200 23074 180000
rect 31942 179200 31998 180000
rect 40866 179200 40922 180000
rect 49790 179200 49846 180000
rect 58714 179200 58770 180000
rect 67638 179200 67694 180000
rect 76562 179200 76618 180000
rect 85486 179200 85542 180000
rect 94410 179200 94466 180000
rect 103334 179200 103390 180000
rect 112258 179200 112314 180000
rect 121182 179200 121238 180000
rect 130106 179200 130162 180000
rect 139030 179200 139086 180000
rect 147954 179200 148010 180000
rect 156878 179200 156934 180000
rect 165802 179200 165858 180000
rect 174726 179200 174782 180000
rect 4986 0 5042 800
rect 13082 0 13138 800
rect 21178 0 21234 800
rect 29274 0 29330 800
rect 37370 0 37426 800
rect 45466 0 45522 800
rect 53562 0 53618 800
rect 61658 0 61714 800
rect 69754 0 69810 800
rect 77850 0 77906 800
rect 85946 0 86002 800
rect 94042 0 94098 800
rect 102138 0 102194 800
rect 110234 0 110290 800
rect 118330 0 118386 800
rect 126426 0 126482 800
rect 134522 0 134578 800
rect 142618 0 142674 800
rect 150714 0 150770 800
rect 158810 0 158866 800
rect 166906 0 166962 800
rect 175002 0 175058 800
<< obsm2 >>
rect 1306 179144 5114 179330
rect 5282 179144 14038 179330
rect 14206 179144 22962 179330
rect 23130 179144 31886 179330
rect 32054 179144 40810 179330
rect 40978 179144 49734 179330
rect 49902 179144 58658 179330
rect 58826 179144 67582 179330
rect 67750 179144 76506 179330
rect 76674 179144 85430 179330
rect 85598 179144 94354 179330
rect 94522 179144 103278 179330
rect 103446 179144 112202 179330
rect 112370 179144 121126 179330
rect 121294 179144 130050 179330
rect 130218 179144 138974 179330
rect 139142 179144 147898 179330
rect 148066 179144 156822 179330
rect 156990 179144 165746 179330
rect 165914 179144 174670 179330
rect 174838 179144 178370 179330
rect 1306 856 178370 179144
rect 1306 800 4930 856
rect 5098 800 13026 856
rect 13194 800 21122 856
rect 21290 800 29218 856
rect 29386 800 37314 856
rect 37482 800 45410 856
rect 45578 800 53506 856
rect 53674 800 61602 856
rect 61770 800 69698 856
rect 69866 800 77794 856
rect 77962 800 85890 856
rect 86058 800 93986 856
rect 94154 800 102082 856
rect 102250 800 110178 856
rect 110346 800 118274 856
rect 118442 800 126370 856
rect 126538 800 134466 856
rect 134634 800 142562 856
rect 142730 800 150658 856
rect 150826 800 158754 856
rect 158922 800 166850 856
rect 167018 800 174946 856
rect 175114 800 178370 856
<< metal3 >>
rect 0 175584 800 175704
rect 179200 175584 180000 175704
rect 0 167424 800 167544
rect 179200 167424 180000 167544
rect 0 159264 800 159384
rect 179200 159264 180000 159384
rect 0 151104 800 151224
rect 179200 151104 180000 151224
rect 0 142944 800 143064
rect 179200 142944 180000 143064
rect 0 134784 800 134904
rect 179200 134784 180000 134904
rect 0 126624 800 126744
rect 179200 126624 180000 126744
rect 0 118464 800 118584
rect 179200 118464 180000 118584
rect 0 110304 800 110424
rect 179200 110304 180000 110424
rect 0 102144 800 102264
rect 179200 102144 180000 102264
rect 0 93984 800 94104
rect 179200 93984 180000 94104
rect 0 85824 800 85944
rect 179200 85824 180000 85944
rect 0 77664 800 77784
rect 179200 77664 180000 77784
rect 0 69504 800 69624
rect 179200 69504 180000 69624
rect 0 61344 800 61464
rect 179200 61344 180000 61464
rect 0 53184 800 53304
rect 179200 53184 180000 53304
rect 0 45024 800 45144
rect 179200 45024 180000 45144
rect 0 36864 800 36984
rect 179200 36864 180000 36984
rect 0 28704 800 28824
rect 179200 28704 180000 28824
rect 0 20544 800 20664
rect 179200 20544 180000 20664
rect 0 12384 800 12504
rect 179200 12384 180000 12504
rect 0 4224 800 4344
rect 179200 4224 180000 4344
<< obsm3 >>
rect 800 175784 179200 177377
rect 880 175504 179120 175784
rect 800 167624 179200 175504
rect 880 167344 179120 167624
rect 800 159464 179200 167344
rect 880 159184 179120 159464
rect 800 151304 179200 159184
rect 880 151024 179120 151304
rect 800 143144 179200 151024
rect 880 142864 179120 143144
rect 800 134984 179200 142864
rect 880 134704 179120 134984
rect 800 126824 179200 134704
rect 880 126544 179120 126824
rect 800 118664 179200 126544
rect 880 118384 179120 118664
rect 800 110504 179200 118384
rect 880 110224 179120 110504
rect 800 102344 179200 110224
rect 880 102064 179120 102344
rect 800 94184 179200 102064
rect 880 93904 179120 94184
rect 800 86024 179200 93904
rect 880 85744 179120 86024
rect 800 77864 179200 85744
rect 880 77584 179120 77864
rect 800 69704 179200 77584
rect 880 69424 179120 69704
rect 800 61544 179200 69424
rect 880 61264 179120 61544
rect 800 53384 179200 61264
rect 880 53104 179120 53384
rect 800 45224 179200 53104
rect 880 44944 179120 45224
rect 800 37064 179200 44944
rect 880 36784 179120 37064
rect 800 28904 179200 36784
rect 880 28624 179120 28904
rect 800 20744 179200 28624
rect 880 20464 179120 20744
rect 800 12584 179200 20464
rect 880 12304 179120 12584
rect 800 4424 179200 12304
rect 880 4144 179120 4424
rect 800 2143 179200 4144
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
<< obsm4 >>
rect 1715 45459 4128 159493
rect 4608 45459 19488 159493
rect 19968 45459 34848 159493
rect 35328 45459 50208 159493
rect 50688 45459 65568 159493
rect 66048 45459 80928 159493
rect 81408 45459 96288 159493
rect 96768 45459 111648 159493
rect 112128 45459 127008 159493
rect 127488 45459 142368 159493
rect 142848 45459 157728 159493
rect 158208 45459 173088 159493
rect 173568 45459 177869 159493
<< labels >>
rlabel metal2 s 4986 0 5042 800 6 hold
port 1 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 iclk
port 2 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 idata
port 3 nsew signal input
rlabel metal3 s 179200 4224 180000 4344 6 ieast[0]
port 4 nsew signal input
rlabel metal3 s 179200 12384 180000 12504 6 ieast[1]
port 5 nsew signal input
rlabel metal3 s 179200 20544 180000 20664 6 ieast[2]
port 6 nsew signal input
rlabel metal3 s 179200 28704 180000 28824 6 ieast[3]
port 7 nsew signal input
rlabel metal3 s 179200 36864 180000 36984 6 ieast[4]
port 8 nsew signal input
rlabel metal3 s 179200 45024 180000 45144 6 ieast[5]
port 9 nsew signal input
rlabel metal3 s 179200 53184 180000 53304 6 ieast[6]
port 10 nsew signal input
rlabel metal3 s 179200 61344 180000 61464 6 ieast[7]
port 11 nsew signal input
rlabel metal3 s 179200 69504 180000 69624 6 ieast[8]
port 12 nsew signal input
rlabel metal3 s 179200 77664 180000 77784 6 ieast[9]
port 13 nsew signal input
rlabel metal2 s 174726 179200 174782 180000 6 inorth[0]
port 14 nsew signal input
rlabel metal2 s 165802 179200 165858 180000 6 inorth[1]
port 15 nsew signal input
rlabel metal2 s 156878 179200 156934 180000 6 inorth[2]
port 16 nsew signal input
rlabel metal2 s 147954 179200 148010 180000 6 inorth[3]
port 17 nsew signal input
rlabel metal2 s 139030 179200 139086 180000 6 inorth[4]
port 18 nsew signal input
rlabel metal2 s 130106 179200 130162 180000 6 inorth[5]
port 19 nsew signal input
rlabel metal2 s 121182 179200 121238 180000 6 inorth[6]
port 20 nsew signal input
rlabel metal2 s 112258 179200 112314 180000 6 inorth[7]
port 21 nsew signal input
rlabel metal2 s 103334 179200 103390 180000 6 inorth[8]
port 22 nsew signal input
rlabel metal2 s 94410 179200 94466 180000 6 inorth[9]
port 23 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 isouth[0]
port 24 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 isouth[1]
port 25 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 isouth[2]
port 26 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 isouth[3]
port 27 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 isouth[4]
port 28 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 isouth[5]
port 29 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 isouth[6]
port 30 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 isouth[7]
port 31 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 isouth[8]
port 32 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 isouth[9]
port 33 nsew signal input
rlabel metal3 s 0 175584 800 175704 6 iwest[0]
port 34 nsew signal input
rlabel metal3 s 0 167424 800 167544 6 iwest[1]
port 35 nsew signal input
rlabel metal3 s 0 159264 800 159384 6 iwest[2]
port 36 nsew signal input
rlabel metal3 s 0 151104 800 151224 6 iwest[3]
port 37 nsew signal input
rlabel metal3 s 0 142944 800 143064 6 iwest[4]
port 38 nsew signal input
rlabel metal3 s 0 134784 800 134904 6 iwest[5]
port 39 nsew signal input
rlabel metal3 s 0 126624 800 126744 6 iwest[6]
port 40 nsew signal input
rlabel metal3 s 0 118464 800 118584 6 iwest[7]
port 41 nsew signal input
rlabel metal3 s 0 110304 800 110424 6 iwest[8]
port 42 nsew signal input
rlabel metal3 s 0 102144 800 102264 6 iwest[9]
port 43 nsew signal input
rlabel metal3 s 179200 167424 180000 167544 6 oclk
port 44 nsew signal output
rlabel metal3 s 179200 175584 180000 175704 6 odata
port 45 nsew signal output
rlabel metal3 s 179200 85824 180000 85944 6 oeast[0]
port 46 nsew signal output
rlabel metal3 s 179200 93984 180000 94104 6 oeast[1]
port 47 nsew signal output
rlabel metal3 s 179200 102144 180000 102264 6 oeast[2]
port 48 nsew signal output
rlabel metal3 s 179200 110304 180000 110424 6 oeast[3]
port 49 nsew signal output
rlabel metal3 s 179200 118464 180000 118584 6 oeast[4]
port 50 nsew signal output
rlabel metal3 s 179200 126624 180000 126744 6 oeast[5]
port 51 nsew signal output
rlabel metal3 s 179200 134784 180000 134904 6 oeast[6]
port 52 nsew signal output
rlabel metal3 s 179200 142944 180000 143064 6 oeast[7]
port 53 nsew signal output
rlabel metal3 s 179200 151104 180000 151224 6 oeast[8]
port 54 nsew signal output
rlabel metal3 s 179200 159264 180000 159384 6 oeast[9]
port 55 nsew signal output
rlabel metal2 s 85486 179200 85542 180000 6 onorth[0]
port 56 nsew signal output
rlabel metal2 s 76562 179200 76618 180000 6 onorth[1]
port 57 nsew signal output
rlabel metal2 s 67638 179200 67694 180000 6 onorth[2]
port 58 nsew signal output
rlabel metal2 s 58714 179200 58770 180000 6 onorth[3]
port 59 nsew signal output
rlabel metal2 s 49790 179200 49846 180000 6 onorth[4]
port 60 nsew signal output
rlabel metal2 s 40866 179200 40922 180000 6 onorth[5]
port 61 nsew signal output
rlabel metal2 s 31942 179200 31998 180000 6 onorth[6]
port 62 nsew signal output
rlabel metal2 s 23018 179200 23074 180000 6 onorth[7]
port 63 nsew signal output
rlabel metal2 s 14094 179200 14150 180000 6 onorth[8]
port 64 nsew signal output
rlabel metal2 s 5170 179200 5226 180000 6 onorth[9]
port 65 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 osouth[0]
port 66 nsew signal output
rlabel metal2 s 110234 0 110290 800 6 osouth[1]
port 67 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 osouth[2]
port 68 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 osouth[3]
port 69 nsew signal output
rlabel metal2 s 134522 0 134578 800 6 osouth[4]
port 70 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 osouth[5]
port 71 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 osouth[6]
port 72 nsew signal output
rlabel metal2 s 158810 0 158866 800 6 osouth[7]
port 73 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 osouth[8]
port 74 nsew signal output
rlabel metal2 s 175002 0 175058 800 6 osouth[9]
port 75 nsew signal output
rlabel metal3 s 0 93984 800 94104 6 owest[0]
port 76 nsew signal output
rlabel metal3 s 0 85824 800 85944 6 owest[1]
port 77 nsew signal output
rlabel metal3 s 0 77664 800 77784 6 owest[2]
port 78 nsew signal output
rlabel metal3 s 0 69504 800 69624 6 owest[3]
port 79 nsew signal output
rlabel metal3 s 0 61344 800 61464 6 owest[4]
port 80 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 owest[5]
port 81 nsew signal output
rlabel metal3 s 0 45024 800 45144 6 owest[6]
port 82 nsew signal output
rlabel metal3 s 0 36864 800 36984 6 owest[7]
port 83 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 owest[8]
port 84 nsew signal output
rlabel metal3 s 0 20544 800 20664 6 owest[9]
port 85 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 reset
port 86 nsew signal input
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 177392 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 177392 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 177392 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 177392 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 177392 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 177392 6 vssd1
port 88 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 38801798
string GDS_FILE /home/alex/chaos_automaton_Summer_2022/openlane/chaos_subarray/runs/22_08_04_13_04/results/signoff/chaos_subarray.magic.gds
string GDS_START 141920
<< end >>

