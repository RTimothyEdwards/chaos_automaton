magic
tech minimum
timestamp 0
<< checkpaint >>
rect 0 0 1 1
<< end >>
